magic
tech gf180mcuC
magscale 1 5
timestamp 1670229454
<< obsm1 >>
rect 10672 2087 149903 106757
<< metal2 >>
rect 4900 299760 5012 300480
rect 13188 299760 13300 300480
rect 21476 299760 21588 300480
rect 38052 299760 38164 300480
rect 46340 299760 46452 300480
rect 54628 299760 54740 300480
rect 71204 299760 71316 300480
rect 79492 299760 79604 300480
rect 87780 299760 87892 300480
rect 104356 299760 104468 300480
rect 112644 299760 112756 300480
rect 120932 299760 121044 300480
rect 137508 299760 137620 300480
rect 145796 299760 145908 300480
rect 154084 299760 154196 300480
rect 170660 299760 170772 300480
rect 178948 299760 179060 300480
rect 187236 299760 187348 300480
rect 203812 299760 203924 300480
rect 212100 299760 212212 300480
rect 220388 299760 220500 300480
rect 236964 299760 237076 300480
rect 245252 299760 245364 300480
rect 253540 299760 253652 300480
rect 270116 299760 270228 300480
rect 278404 299760 278516 300480
rect 286692 299760 286804 300480
rect 11900 -480 12012 240
rect 12460 -480 12572 240
rect 13020 -480 13132 240
rect 13580 -480 13692 240
rect 14140 -480 14252 240
rect 14700 -480 14812 240
rect 15260 -480 15372 240
rect 15820 -480 15932 240
rect 16380 -480 16492 240
rect 16940 -480 17052 240
rect 17500 -480 17612 240
rect 18060 -480 18172 240
rect 18620 -480 18732 240
rect 19180 -480 19292 240
rect 19740 -480 19852 240
rect 20300 -480 20412 240
rect 20860 -480 20972 240
rect 21420 -480 21532 240
rect 21980 -480 22092 240
rect 22540 -480 22652 240
rect 23100 -480 23212 240
rect 23660 -480 23772 240
rect 24220 -480 24332 240
rect 24780 -480 24892 240
rect 25340 -480 25452 240
rect 25900 -480 26012 240
rect 26460 -480 26572 240
rect 27020 -480 27132 240
rect 27580 -480 27692 240
rect 28140 -480 28252 240
rect 28700 -480 28812 240
rect 29260 -480 29372 240
rect 29820 -480 29932 240
rect 30380 -480 30492 240
rect 30940 -480 31052 240
rect 31500 -480 31612 240
rect 32060 -480 32172 240
rect 32620 -480 32732 240
rect 33180 -480 33292 240
rect 33740 -480 33852 240
rect 34300 -480 34412 240
rect 34860 -480 34972 240
rect 35420 -480 35532 240
rect 35980 -480 36092 240
rect 36540 -480 36652 240
rect 37100 -480 37212 240
rect 37660 -480 37772 240
rect 38220 -480 38332 240
rect 38780 -480 38892 240
rect 39340 -480 39452 240
rect 39900 -480 40012 240
rect 40460 -480 40572 240
rect 41020 -480 41132 240
rect 41580 -480 41692 240
rect 42140 -480 42252 240
rect 42700 -480 42812 240
rect 43260 -480 43372 240
rect 43820 -480 43932 240
rect 44380 -480 44492 240
rect 44940 -480 45052 240
rect 45500 -480 45612 240
rect 46060 -480 46172 240
rect 46620 -480 46732 240
rect 47180 -480 47292 240
rect 47740 -480 47852 240
rect 48300 -480 48412 240
rect 48860 -480 48972 240
rect 49420 -480 49532 240
rect 49980 -480 50092 240
rect 50540 -480 50652 240
rect 51100 -480 51212 240
rect 51660 -480 51772 240
rect 52220 -480 52332 240
rect 52780 -480 52892 240
rect 53340 -480 53452 240
rect 53900 -480 54012 240
rect 54460 -480 54572 240
rect 55020 -480 55132 240
rect 55580 -480 55692 240
rect 56140 -480 56252 240
rect 56700 -480 56812 240
rect 57260 -480 57372 240
rect 57820 -480 57932 240
rect 58380 -480 58492 240
rect 58940 -480 59052 240
rect 59500 -480 59612 240
rect 60060 -480 60172 240
rect 60620 -480 60732 240
rect 61180 -480 61292 240
rect 61740 -480 61852 240
rect 62300 -480 62412 240
rect 62860 -480 62972 240
rect 63420 -480 63532 240
rect 63980 -480 64092 240
rect 64540 -480 64652 240
rect 65100 -480 65212 240
rect 65660 -480 65772 240
rect 66220 -480 66332 240
rect 66780 -480 66892 240
rect 67340 -480 67452 240
rect 67900 -480 68012 240
rect 68460 -480 68572 240
rect 69020 -480 69132 240
rect 69580 -480 69692 240
rect 70140 -480 70252 240
rect 70700 -480 70812 240
rect 71260 -480 71372 240
rect 71820 -480 71932 240
rect 72380 -480 72492 240
rect 72940 -480 73052 240
rect 73500 -480 73612 240
rect 74060 -480 74172 240
rect 74620 -480 74732 240
rect 75180 -480 75292 240
rect 75740 -480 75852 240
rect 76300 -480 76412 240
rect 76860 -480 76972 240
rect 77420 -480 77532 240
rect 77980 -480 78092 240
rect 78540 -480 78652 240
rect 79100 -480 79212 240
rect 79660 -480 79772 240
rect 80220 -480 80332 240
rect 80780 -480 80892 240
rect 81340 -480 81452 240
rect 81900 -480 82012 240
rect 82460 -480 82572 240
rect 83020 -480 83132 240
rect 83580 -480 83692 240
rect 84140 -480 84252 240
rect 84700 -480 84812 240
rect 85260 -480 85372 240
rect 85820 -480 85932 240
rect 86380 -480 86492 240
rect 86940 -480 87052 240
rect 87500 -480 87612 240
rect 88060 -480 88172 240
rect 88620 -480 88732 240
rect 89180 -480 89292 240
rect 89740 -480 89852 240
rect 90300 -480 90412 240
rect 90860 -480 90972 240
rect 91420 -480 91532 240
rect 91980 -480 92092 240
rect 92540 -480 92652 240
rect 93100 -480 93212 240
rect 93660 -480 93772 240
rect 94220 -480 94332 240
rect 94780 -480 94892 240
rect 95340 -480 95452 240
rect 95900 -480 96012 240
rect 96460 -480 96572 240
rect 97020 -480 97132 240
rect 97580 -480 97692 240
rect 98140 -480 98252 240
rect 98700 -480 98812 240
rect 99260 -480 99372 240
rect 99820 -480 99932 240
rect 100380 -480 100492 240
rect 100940 -480 101052 240
rect 101500 -480 101612 240
rect 102060 -480 102172 240
rect 102620 -480 102732 240
rect 103180 -480 103292 240
rect 103740 -480 103852 240
rect 104300 -480 104412 240
rect 104860 -480 104972 240
rect 105420 -480 105532 240
rect 105980 -480 106092 240
rect 106540 -480 106652 240
rect 107100 -480 107212 240
rect 107660 -480 107772 240
rect 108220 -480 108332 240
rect 108780 -480 108892 240
rect 109340 -480 109452 240
rect 109900 -480 110012 240
rect 110460 -480 110572 240
rect 111020 -480 111132 240
rect 111580 -480 111692 240
rect 112140 -480 112252 240
rect 112700 -480 112812 240
rect 113260 -480 113372 240
rect 113820 -480 113932 240
rect 114380 -480 114492 240
rect 114940 -480 115052 240
rect 115500 -480 115612 240
rect 116060 -480 116172 240
rect 116620 -480 116732 240
rect 117180 -480 117292 240
rect 117740 -480 117852 240
rect 118300 -480 118412 240
rect 118860 -480 118972 240
rect 119420 -480 119532 240
rect 119980 -480 120092 240
rect 120540 -480 120652 240
rect 121100 -480 121212 240
rect 121660 -480 121772 240
rect 122220 -480 122332 240
rect 122780 -480 122892 240
rect 123340 -480 123452 240
rect 123900 -480 124012 240
rect 124460 -480 124572 240
rect 125020 -480 125132 240
rect 125580 -480 125692 240
rect 126140 -480 126252 240
rect 126700 -480 126812 240
rect 127260 -480 127372 240
rect 127820 -480 127932 240
rect 128380 -480 128492 240
rect 128940 -480 129052 240
rect 129500 -480 129612 240
rect 130060 -480 130172 240
rect 130620 -480 130732 240
rect 131180 -480 131292 240
rect 131740 -480 131852 240
rect 132300 -480 132412 240
rect 132860 -480 132972 240
rect 133420 -480 133532 240
rect 133980 -480 134092 240
rect 134540 -480 134652 240
rect 135100 -480 135212 240
rect 135660 -480 135772 240
rect 136220 -480 136332 240
rect 136780 -480 136892 240
rect 137340 -480 137452 240
rect 137900 -480 138012 240
rect 138460 -480 138572 240
rect 139020 -480 139132 240
rect 139580 -480 139692 240
rect 140140 -480 140252 240
rect 140700 -480 140812 240
rect 141260 -480 141372 240
rect 141820 -480 141932 240
rect 142380 -480 142492 240
rect 142940 -480 143052 240
rect 143500 -480 143612 240
rect 144060 -480 144172 240
rect 144620 -480 144732 240
rect 145180 -480 145292 240
rect 145740 -480 145852 240
rect 146300 -480 146412 240
rect 146860 -480 146972 240
rect 147420 -480 147532 240
rect 147980 -480 148092 240
rect 148540 -480 148652 240
rect 149100 -480 149212 240
rect 149660 -480 149772 240
rect 150220 -480 150332 240
rect 150780 -480 150892 240
rect 151340 -480 151452 240
rect 151900 -480 152012 240
rect 152460 -480 152572 240
rect 153020 -480 153132 240
rect 153580 -480 153692 240
rect 154140 -480 154252 240
rect 154700 -480 154812 240
rect 155260 -480 155372 240
rect 155820 -480 155932 240
rect 156380 -480 156492 240
rect 156940 -480 157052 240
rect 157500 -480 157612 240
rect 158060 -480 158172 240
rect 158620 -480 158732 240
rect 159180 -480 159292 240
rect 159740 -480 159852 240
rect 160300 -480 160412 240
rect 160860 -480 160972 240
rect 161420 -480 161532 240
rect 161980 -480 162092 240
rect 162540 -480 162652 240
rect 163100 -480 163212 240
rect 163660 -480 163772 240
rect 164220 -480 164332 240
rect 164780 -480 164892 240
rect 165340 -480 165452 240
rect 165900 -480 166012 240
rect 166460 -480 166572 240
rect 167020 -480 167132 240
rect 167580 -480 167692 240
rect 168140 -480 168252 240
rect 168700 -480 168812 240
rect 169260 -480 169372 240
rect 169820 -480 169932 240
rect 170380 -480 170492 240
rect 170940 -480 171052 240
rect 171500 -480 171612 240
rect 172060 -480 172172 240
rect 172620 -480 172732 240
rect 173180 -480 173292 240
rect 173740 -480 173852 240
rect 174300 -480 174412 240
rect 174860 -480 174972 240
rect 175420 -480 175532 240
rect 175980 -480 176092 240
rect 176540 -480 176652 240
rect 177100 -480 177212 240
rect 177660 -480 177772 240
rect 178220 -480 178332 240
rect 286300 -480 286412 240
rect 286860 -480 286972 240
rect 287420 -480 287532 240
rect 287980 -480 288092 240
<< obsm2 >>
rect 14 299730 4870 299810
rect 5042 299730 13158 299810
rect 13330 299730 21446 299810
rect 21618 299730 38022 299810
rect 38194 299730 46310 299810
rect 46482 299730 54598 299810
rect 54770 299730 71174 299810
rect 71346 299730 79462 299810
rect 79634 299730 87750 299810
rect 87922 299730 104326 299810
rect 104498 299730 112614 299810
rect 112786 299730 120902 299810
rect 121074 299730 137478 299810
rect 137650 299730 145766 299810
rect 145938 299730 154054 299810
rect 154226 299730 170630 299810
rect 170802 299730 178918 299810
rect 179090 299730 187206 299810
rect 187378 299730 203782 299810
rect 203954 299730 212070 299810
rect 212242 299730 220358 299810
rect 220530 299730 236934 299810
rect 237106 299730 245222 299810
rect 245394 299730 253510 299810
rect 253682 299730 270086 299810
rect 270258 299730 278374 299810
rect 278546 299730 286662 299810
rect 286834 299730 299586 299810
rect 14 270 299586 299730
rect 14 9 11870 270
rect 12042 9 12430 270
rect 12602 9 12990 270
rect 13162 9 13550 270
rect 13722 9 14110 270
rect 14282 9 14670 270
rect 14842 9 15230 270
rect 15402 9 15790 270
rect 15962 9 16350 270
rect 16522 9 16910 270
rect 17082 9 17470 270
rect 17642 9 18030 270
rect 18202 9 18590 270
rect 18762 9 19150 270
rect 19322 9 19710 270
rect 19882 9 20270 270
rect 20442 9 20830 270
rect 21002 9 21390 270
rect 21562 9 21950 270
rect 22122 9 22510 270
rect 22682 9 23070 270
rect 23242 9 23630 270
rect 23802 9 24190 270
rect 24362 9 24750 270
rect 24922 9 25310 270
rect 25482 9 25870 270
rect 26042 9 26430 270
rect 26602 9 26990 270
rect 27162 9 27550 270
rect 27722 9 28110 270
rect 28282 9 28670 270
rect 28842 9 29230 270
rect 29402 9 29790 270
rect 29962 9 30350 270
rect 30522 9 30910 270
rect 31082 9 31470 270
rect 31642 9 32030 270
rect 32202 9 32590 270
rect 32762 9 33150 270
rect 33322 9 33710 270
rect 33882 9 34270 270
rect 34442 9 34830 270
rect 35002 9 35390 270
rect 35562 9 35950 270
rect 36122 9 36510 270
rect 36682 9 37070 270
rect 37242 9 37630 270
rect 37802 9 38190 270
rect 38362 9 38750 270
rect 38922 9 39310 270
rect 39482 9 39870 270
rect 40042 9 40430 270
rect 40602 9 40990 270
rect 41162 9 41550 270
rect 41722 9 42110 270
rect 42282 9 42670 270
rect 42842 9 43230 270
rect 43402 9 43790 270
rect 43962 9 44350 270
rect 44522 9 44910 270
rect 45082 9 45470 270
rect 45642 9 46030 270
rect 46202 9 46590 270
rect 46762 9 47150 270
rect 47322 9 47710 270
rect 47882 9 48270 270
rect 48442 9 48830 270
rect 49002 9 49390 270
rect 49562 9 49950 270
rect 50122 9 50510 270
rect 50682 9 51070 270
rect 51242 9 51630 270
rect 51802 9 52190 270
rect 52362 9 52750 270
rect 52922 9 53310 270
rect 53482 9 53870 270
rect 54042 9 54430 270
rect 54602 9 54990 270
rect 55162 9 55550 270
rect 55722 9 56110 270
rect 56282 9 56670 270
rect 56842 9 57230 270
rect 57402 9 57790 270
rect 57962 9 58350 270
rect 58522 9 58910 270
rect 59082 9 59470 270
rect 59642 9 60030 270
rect 60202 9 60590 270
rect 60762 9 61150 270
rect 61322 9 61710 270
rect 61882 9 62270 270
rect 62442 9 62830 270
rect 63002 9 63390 270
rect 63562 9 63950 270
rect 64122 9 64510 270
rect 64682 9 65070 270
rect 65242 9 65630 270
rect 65802 9 66190 270
rect 66362 9 66750 270
rect 66922 9 67310 270
rect 67482 9 67870 270
rect 68042 9 68430 270
rect 68602 9 68990 270
rect 69162 9 69550 270
rect 69722 9 70110 270
rect 70282 9 70670 270
rect 70842 9 71230 270
rect 71402 9 71790 270
rect 71962 9 72350 270
rect 72522 9 72910 270
rect 73082 9 73470 270
rect 73642 9 74030 270
rect 74202 9 74590 270
rect 74762 9 75150 270
rect 75322 9 75710 270
rect 75882 9 76270 270
rect 76442 9 76830 270
rect 77002 9 77390 270
rect 77562 9 77950 270
rect 78122 9 78510 270
rect 78682 9 79070 270
rect 79242 9 79630 270
rect 79802 9 80190 270
rect 80362 9 80750 270
rect 80922 9 81310 270
rect 81482 9 81870 270
rect 82042 9 82430 270
rect 82602 9 82990 270
rect 83162 9 83550 270
rect 83722 9 84110 270
rect 84282 9 84670 270
rect 84842 9 85230 270
rect 85402 9 85790 270
rect 85962 9 86350 270
rect 86522 9 86910 270
rect 87082 9 87470 270
rect 87642 9 88030 270
rect 88202 9 88590 270
rect 88762 9 89150 270
rect 89322 9 89710 270
rect 89882 9 90270 270
rect 90442 9 90830 270
rect 91002 9 91390 270
rect 91562 9 91950 270
rect 92122 9 92510 270
rect 92682 9 93070 270
rect 93242 9 93630 270
rect 93802 9 94190 270
rect 94362 9 94750 270
rect 94922 9 95310 270
rect 95482 9 95870 270
rect 96042 9 96430 270
rect 96602 9 96990 270
rect 97162 9 97550 270
rect 97722 9 98110 270
rect 98282 9 98670 270
rect 98842 9 99230 270
rect 99402 9 99790 270
rect 99962 9 100350 270
rect 100522 9 100910 270
rect 101082 9 101470 270
rect 101642 9 102030 270
rect 102202 9 102590 270
rect 102762 9 103150 270
rect 103322 9 103710 270
rect 103882 9 104270 270
rect 104442 9 104830 270
rect 105002 9 105390 270
rect 105562 9 105950 270
rect 106122 9 106510 270
rect 106682 9 107070 270
rect 107242 9 107630 270
rect 107802 9 108190 270
rect 108362 9 108750 270
rect 108922 9 109310 270
rect 109482 9 109870 270
rect 110042 9 110430 270
rect 110602 9 110990 270
rect 111162 9 111550 270
rect 111722 9 112110 270
rect 112282 9 112670 270
rect 112842 9 113230 270
rect 113402 9 113790 270
rect 113962 9 114350 270
rect 114522 9 114910 270
rect 115082 9 115470 270
rect 115642 9 116030 270
rect 116202 9 116590 270
rect 116762 9 117150 270
rect 117322 9 117710 270
rect 117882 9 118270 270
rect 118442 9 118830 270
rect 119002 9 119390 270
rect 119562 9 119950 270
rect 120122 9 120510 270
rect 120682 9 121070 270
rect 121242 9 121630 270
rect 121802 9 122190 270
rect 122362 9 122750 270
rect 122922 9 123310 270
rect 123482 9 123870 270
rect 124042 9 124430 270
rect 124602 9 124990 270
rect 125162 9 125550 270
rect 125722 9 126110 270
rect 126282 9 126670 270
rect 126842 9 127230 270
rect 127402 9 127790 270
rect 127962 9 128350 270
rect 128522 9 128910 270
rect 129082 9 129470 270
rect 129642 9 130030 270
rect 130202 9 130590 270
rect 130762 9 131150 270
rect 131322 9 131710 270
rect 131882 9 132270 270
rect 132442 9 132830 270
rect 133002 9 133390 270
rect 133562 9 133950 270
rect 134122 9 134510 270
rect 134682 9 135070 270
rect 135242 9 135630 270
rect 135802 9 136190 270
rect 136362 9 136750 270
rect 136922 9 137310 270
rect 137482 9 137870 270
rect 138042 9 138430 270
rect 138602 9 138990 270
rect 139162 9 139550 270
rect 139722 9 140110 270
rect 140282 9 140670 270
rect 140842 9 141230 270
rect 141402 9 141790 270
rect 141962 9 142350 270
rect 142522 9 142910 270
rect 143082 9 143470 270
rect 143642 9 144030 270
rect 144202 9 144590 270
rect 144762 9 145150 270
rect 145322 9 145710 270
rect 145882 9 146270 270
rect 146442 9 146830 270
rect 147002 9 147390 270
rect 147562 9 147950 270
rect 148122 9 148510 270
rect 148682 9 149070 270
rect 149242 9 149630 270
rect 149802 9 150190 270
rect 150362 9 150750 270
rect 150922 9 151310 270
rect 151482 9 151870 270
rect 152042 9 152430 270
rect 152602 9 152990 270
rect 153162 9 153550 270
rect 153722 9 154110 270
rect 154282 9 154670 270
rect 154842 9 155230 270
rect 155402 9 155790 270
rect 155962 9 156350 270
rect 156522 9 156910 270
rect 157082 9 157470 270
rect 157642 9 158030 270
rect 158202 9 158590 270
rect 158762 9 159150 270
rect 159322 9 159710 270
rect 159882 9 160270 270
rect 160442 9 160830 270
rect 161002 9 161390 270
rect 161562 9 161950 270
rect 162122 9 162510 270
rect 162682 9 163070 270
rect 163242 9 163630 270
rect 163802 9 164190 270
rect 164362 9 164750 270
rect 164922 9 165310 270
rect 165482 9 165870 270
rect 166042 9 166430 270
rect 166602 9 166990 270
rect 167162 9 167550 270
rect 167722 9 168110 270
rect 168282 9 168670 270
rect 168842 9 169230 270
rect 169402 9 169790 270
rect 169962 9 170350 270
rect 170522 9 170910 270
rect 171082 9 171470 270
rect 171642 9 172030 270
rect 172202 9 172590 270
rect 172762 9 173150 270
rect 173322 9 173710 270
rect 173882 9 174270 270
rect 174442 9 174830 270
rect 175002 9 175390 270
rect 175562 9 175950 270
rect 176122 9 176510 270
rect 176682 9 177070 270
rect 177242 9 177630 270
rect 177802 9 178190 270
rect 178362 9 286270 270
rect 286442 9 286830 270
rect 287002 9 287390 270
rect 287562 9 287950 270
rect 288122 9 299586 270
<< metal3 >>
rect 299760 296996 300480 297108
rect -480 291284 240 291396
rect 299760 291340 300480 291452
rect -480 285740 240 285852
rect 299760 285684 300480 285796
rect -480 280196 240 280308
rect 299760 274372 300480 274484
rect -480 269108 240 269220
rect 299760 268716 300480 268828
rect -480 263564 240 263676
rect 299760 263060 300480 263172
rect -480 258020 240 258132
rect 299760 251748 300480 251860
rect -480 246932 240 247044
rect 299760 246092 300480 246204
rect -480 241388 240 241500
rect 299760 240436 300480 240548
rect -480 235844 240 235956
rect 299760 229124 300480 229236
rect -480 224756 240 224868
rect 299760 223468 300480 223580
rect -480 219212 240 219324
rect 299760 217812 300480 217924
rect -480 213668 240 213780
rect 299760 206500 300480 206612
rect -480 202580 240 202692
rect 299760 200844 300480 200956
rect -480 197036 240 197148
rect 299760 195188 300480 195300
rect -480 191492 240 191604
rect 299760 183876 300480 183988
rect -480 180404 240 180516
rect 299760 178220 300480 178332
rect -480 174860 240 174972
rect 299760 172564 300480 172676
rect -480 169316 240 169428
rect 299760 161252 300480 161364
rect -480 158228 240 158340
rect 299760 155596 300480 155708
rect -480 152684 240 152796
rect 299760 149940 300480 150052
rect -480 147140 240 147252
rect 299760 138628 300480 138740
rect -480 136052 240 136164
rect 299760 132972 300480 133084
rect -480 130508 240 130620
rect 299760 127316 300480 127428
rect -480 124964 240 125076
rect 299760 116004 300480 116116
rect -480 113876 240 113988
rect 299760 110348 300480 110460
rect -480 108332 240 108444
rect 299760 104692 300480 104804
rect -480 102788 240 102900
rect 299760 99036 300480 99148
rect 299760 93380 300480 93492
rect -480 91700 240 91812
rect 299760 87724 300480 87836
rect -480 86156 240 86268
rect 299760 82068 300480 82180
rect -480 80612 240 80724
rect 299760 76412 300480 76524
rect 299760 70756 300480 70868
rect -480 69524 240 69636
rect 299760 65100 300480 65212
rect -480 63980 240 64092
rect 299760 59444 300480 59556
rect -480 58436 240 58548
rect 299760 53788 300480 53900
rect 299760 48132 300480 48244
rect -480 47348 240 47460
rect 299760 42476 300480 42588
rect -480 41804 240 41916
rect 299760 36820 300480 36932
rect -480 36260 240 36372
rect 299760 31164 300480 31276
rect -480 30716 240 30828
rect 299760 25508 300480 25620
rect -480 25172 240 25284
rect 299760 19852 300480 19964
rect -480 19628 240 19740
rect -480 14084 240 14196
rect 299760 14196 300480 14308
rect -480 8540 240 8652
rect 299760 8540 300480 8652
rect -480 2996 240 3108
rect 299760 2884 300480 2996
<< obsm3 >>
rect 9 297138 299810 297906
rect 9 296966 299730 297138
rect 9 291482 299810 296966
rect 9 291426 299730 291482
rect 270 291310 299730 291426
rect 270 291254 299810 291310
rect 9 285882 299810 291254
rect 270 285826 299810 285882
rect 270 285710 299730 285826
rect 9 285654 299730 285710
rect 9 280338 299810 285654
rect 270 280166 299810 280338
rect 9 274514 299810 280166
rect 9 274342 299730 274514
rect 9 269250 299810 274342
rect 270 269078 299810 269250
rect 9 268858 299810 269078
rect 9 268686 299730 268858
rect 9 263706 299810 268686
rect 270 263534 299810 263706
rect 9 263202 299810 263534
rect 9 263030 299730 263202
rect 9 258162 299810 263030
rect 270 257990 299810 258162
rect 9 251890 299810 257990
rect 9 251718 299730 251890
rect 9 247074 299810 251718
rect 270 246902 299810 247074
rect 9 246234 299810 246902
rect 9 246062 299730 246234
rect 9 241530 299810 246062
rect 270 241358 299810 241530
rect 9 240578 299810 241358
rect 9 240406 299730 240578
rect 9 235986 299810 240406
rect 270 235814 299810 235986
rect 9 229266 299810 235814
rect 9 229094 299730 229266
rect 9 224898 299810 229094
rect 270 224726 299810 224898
rect 9 223610 299810 224726
rect 9 223438 299730 223610
rect 9 219354 299810 223438
rect 270 219182 299810 219354
rect 9 217954 299810 219182
rect 9 217782 299730 217954
rect 9 213810 299810 217782
rect 270 213638 299810 213810
rect 9 206642 299810 213638
rect 9 206470 299730 206642
rect 9 202722 299810 206470
rect 270 202550 299810 202722
rect 9 200986 299810 202550
rect 9 200814 299730 200986
rect 9 197178 299810 200814
rect 270 197006 299810 197178
rect 9 195330 299810 197006
rect 9 195158 299730 195330
rect 9 191634 299810 195158
rect 270 191462 299810 191634
rect 9 184018 299810 191462
rect 9 183846 299730 184018
rect 9 180546 299810 183846
rect 270 180374 299810 180546
rect 9 178362 299810 180374
rect 9 178190 299730 178362
rect 9 175002 299810 178190
rect 270 174830 299810 175002
rect 9 172706 299810 174830
rect 9 172534 299730 172706
rect 9 169458 299810 172534
rect 270 169286 299810 169458
rect 9 161394 299810 169286
rect 9 161222 299730 161394
rect 9 158370 299810 161222
rect 270 158198 299810 158370
rect 9 155738 299810 158198
rect 9 155566 299730 155738
rect 9 152826 299810 155566
rect 270 152654 299810 152826
rect 9 150082 299810 152654
rect 9 149910 299730 150082
rect 9 147282 299810 149910
rect 270 147110 299810 147282
rect 9 138770 299810 147110
rect 9 138598 299730 138770
rect 9 136194 299810 138598
rect 270 136022 299810 136194
rect 9 133114 299810 136022
rect 9 132942 299730 133114
rect 9 130650 299810 132942
rect 270 130478 299810 130650
rect 9 127458 299810 130478
rect 9 127286 299730 127458
rect 9 125106 299810 127286
rect 270 124934 299810 125106
rect 9 116146 299810 124934
rect 9 115974 299730 116146
rect 9 114018 299810 115974
rect 270 113846 299810 114018
rect 9 110490 299810 113846
rect 9 110318 299730 110490
rect 9 108474 299810 110318
rect 270 108302 299810 108474
rect 9 104834 299810 108302
rect 9 104662 299730 104834
rect 9 102930 299810 104662
rect 270 102758 299810 102930
rect 9 99178 299810 102758
rect 9 99006 299730 99178
rect 9 93522 299810 99006
rect 9 93350 299730 93522
rect 9 91842 299810 93350
rect 270 91670 299810 91842
rect 9 87866 299810 91670
rect 9 87694 299730 87866
rect 9 86298 299810 87694
rect 270 86126 299810 86298
rect 9 82210 299810 86126
rect 9 82038 299730 82210
rect 9 80754 299810 82038
rect 270 80582 299810 80754
rect 9 76554 299810 80582
rect 9 76382 299730 76554
rect 9 70898 299810 76382
rect 9 70726 299730 70898
rect 9 69666 299810 70726
rect 270 69494 299810 69666
rect 9 65242 299810 69494
rect 9 65070 299730 65242
rect 9 64122 299810 65070
rect 270 63950 299810 64122
rect 9 59586 299810 63950
rect 9 59414 299730 59586
rect 9 58578 299810 59414
rect 270 58406 299810 58578
rect 9 53930 299810 58406
rect 9 53758 299730 53930
rect 9 48274 299810 53758
rect 9 48102 299730 48274
rect 9 47490 299810 48102
rect 270 47318 299810 47490
rect 9 42618 299810 47318
rect 9 42446 299730 42618
rect 9 41946 299810 42446
rect 270 41774 299810 41946
rect 9 36962 299810 41774
rect 9 36790 299730 36962
rect 9 36402 299810 36790
rect 270 36230 299810 36402
rect 9 31306 299810 36230
rect 9 31134 299730 31306
rect 9 30858 299810 31134
rect 270 30686 299810 30858
rect 9 25650 299810 30686
rect 9 25478 299730 25650
rect 9 25314 299810 25478
rect 270 25142 299810 25314
rect 9 19994 299810 25142
rect 9 19822 299730 19994
rect 9 19770 299810 19822
rect 270 19598 299810 19770
rect 9 14338 299810 19598
rect 9 14226 299730 14338
rect 270 14166 299730 14226
rect 270 14054 299810 14166
rect 9 8682 299810 14054
rect 270 8510 299730 8682
rect 9 3138 299810 8510
rect 270 3026 299810 3138
rect 270 2966 299730 3026
rect 9 2854 299730 2966
rect 9 14 299810 2854
<< metal4 >>
rect -3283 -2387 -2973 302267
rect -2803 -1907 -2493 301787
rect -2323 -1427 -2013 301307
rect -1843 -947 -1533 300827
rect -1363 -467 -1053 300347
rect -883 13 -573 299867
rect 1017 -2387 1327 302267
rect 2877 -2387 3187 302267
rect 4737 -2387 5047 302267
rect 6597 -2387 6907 302267
rect 8457 -2387 8767 302267
rect 10317 -2387 10627 302267
rect 19017 -2387 19327 302267
rect 20877 -2387 21187 302267
rect 22737 -2387 23047 302267
rect 24597 -2387 24907 302267
rect 26457 94967 26767 302267
rect 28317 94967 28627 302267
rect 37017 94967 37327 302267
rect 38877 94967 39187 302267
rect 40737 94967 41047 302267
rect 42597 94967 42907 302267
rect 44457 94967 44767 302267
rect 26457 -2387 26767 82289
rect 28317 -2387 28627 82289
rect 37017 -2387 37327 82289
rect 38877 -2387 39187 82289
rect 40737 -2387 41047 82289
rect 42597 59415 42907 82289
rect 44457 59415 44767 82289
rect 46317 59415 46627 302267
rect 55017 59415 55327 302267
rect 56877 59415 57187 302267
rect 58737 59415 59047 302267
rect 42597 -2387 42907 51721
rect 44457 -2387 44767 51721
rect 46317 -2387 46627 51721
rect 55017 -2387 55327 51721
rect 56877 -2387 57187 51721
rect 58737 -2387 59047 51721
rect 60597 -2387 60907 302267
rect 62457 -2387 62767 302267
rect 64317 -2387 64627 302267
rect 73017 -2387 73327 302267
rect 74877 -2387 75187 302267
rect 76737 -2387 77047 302267
rect 78597 -2387 78907 302267
rect 80457 -2387 80767 302267
rect 82317 -2387 82627 302267
rect 91017 -2387 91327 302267
rect 92877 -2387 93187 302267
rect 94737 -2387 95047 302267
rect 96597 -2387 96907 302267
rect 98457 -2387 98767 302267
rect 100317 -2387 100627 302267
rect 109017 -2387 109327 302267
rect 110877 -2387 111187 302267
rect 112737 -2387 113047 302267
rect 114597 -2387 114907 302267
rect 116457 -2387 116767 302267
rect 118317 -2387 118627 302267
rect 127017 -2387 127327 302267
rect 128877 -2387 129187 302267
rect 130737 -2387 131047 302267
rect 132597 -2387 132907 302267
rect 134457 -2387 134767 302267
rect 136317 -2387 136627 302267
rect 145017 -2387 145327 302267
rect 146877 -2387 147187 302267
rect 148737 -2387 149047 302267
rect 150597 -2387 150907 302267
rect 152457 -2387 152767 302267
rect 154317 -2387 154627 302267
rect 163017 -2387 163327 302267
rect 164877 -2387 165187 302267
rect 166737 -2387 167047 302267
rect 168597 -2387 168907 302267
rect 170457 -2387 170767 302267
rect 172317 -2387 172627 302267
rect 181017 -2387 181327 302267
rect 182877 -2387 183187 302267
rect 184737 -2387 185047 302267
rect 186597 -2387 186907 302267
rect 188457 -2387 188767 302267
rect 190317 -2387 190627 302267
rect 199017 -2387 199327 302267
rect 200877 -2387 201187 302267
rect 202737 -2387 203047 302267
rect 204597 -2387 204907 302267
rect 206457 -2387 206767 302267
rect 208317 -2387 208627 302267
rect 217017 -2387 217327 302267
rect 218877 -2387 219187 302267
rect 220737 -2387 221047 302267
rect 222597 -2387 222907 302267
rect 224457 -2387 224767 302267
rect 226317 -2387 226627 302267
rect 235017 -2387 235327 302267
rect 236877 -2387 237187 302267
rect 238737 -2387 239047 302267
rect 240597 -2387 240907 302267
rect 242457 -2387 242767 302267
rect 244317 -2387 244627 302267
rect 253017 -2387 253327 302267
rect 254877 -2387 255187 302267
rect 256737 -2387 257047 302267
rect 258597 -2387 258907 302267
rect 260457 -2387 260767 302267
rect 262317 -2387 262627 302267
rect 271017 -2387 271327 302267
rect 272877 -2387 273187 302267
rect 274737 -2387 275047 302267
rect 276597 -2387 276907 302267
rect 278457 -2387 278767 302267
rect 280317 -2387 280627 302267
rect 289017 -2387 289327 302267
rect 290877 -2387 291187 302267
rect 292737 -2387 293047 302267
rect 294597 -2387 294907 302267
rect 296457 -2387 296767 302267
rect 298317 -2387 298627 302267
rect 300565 13 300875 299867
rect 301045 -467 301355 300347
rect 301525 -947 301835 300827
rect 302005 -1427 302315 301307
rect 302485 -1907 302795 301787
rect 302965 -2387 303275 302267
<< obsm4 >>
rect 11438 9 18987 297799
rect 19357 9 20847 297799
rect 21217 9 22707 297799
rect 23077 9 24567 297799
rect 24937 94937 26427 297799
rect 26797 94937 28287 297799
rect 28657 94937 36987 297799
rect 37357 94937 38847 297799
rect 39217 94937 40707 297799
rect 41077 94937 42567 297799
rect 42937 94937 44427 297799
rect 44797 94937 46287 297799
rect 24937 82319 46287 94937
rect 24937 9 26427 82319
rect 26797 9 28287 82319
rect 28657 9 36987 82319
rect 37357 9 38847 82319
rect 39217 9 40707 82319
rect 41077 59385 42567 82319
rect 42937 59385 44427 82319
rect 44797 59385 46287 82319
rect 46657 59385 54987 297799
rect 55357 59385 56847 297799
rect 57217 59385 58707 297799
rect 59077 59385 60567 297799
rect 41077 51751 60567 59385
rect 41077 9 42567 51751
rect 42937 9 44427 51751
rect 44797 9 46287 51751
rect 46657 9 54987 51751
rect 55357 9 56847 51751
rect 57217 9 58707 51751
rect 59077 9 60567 51751
rect 60937 9 62427 297799
rect 62797 9 64287 297799
rect 64657 9 72987 297799
rect 73357 9 74847 297799
rect 75217 9 76707 297799
rect 77077 9 78567 297799
rect 78937 9 80427 297799
rect 80797 9 82287 297799
rect 82657 9 90987 297799
rect 91357 9 92847 297799
rect 93217 9 94707 297799
rect 95077 9 96567 297799
rect 96937 9 98427 297799
rect 98797 9 100287 297799
rect 100657 9 108987 297799
rect 109357 9 110847 297799
rect 111217 9 112707 297799
rect 113077 9 114567 297799
rect 114937 9 116427 297799
rect 116797 9 118287 297799
rect 118657 9 126987 297799
rect 127357 9 128847 297799
rect 129217 9 130707 297799
rect 131077 9 132567 297799
rect 132937 9 134427 297799
rect 134797 9 136287 297799
rect 136657 9 142058 297799
<< metal5 >>
rect -3283 301957 303275 302267
rect -2803 301477 302795 301787
rect -2323 300997 302315 301307
rect -1843 300517 301835 300827
rect -1363 300037 301355 300347
rect -883 299557 300875 299867
rect -3283 297353 303275 297663
rect -3283 295493 303275 295803
rect -3283 293633 303275 293943
rect -3283 291773 303275 292083
rect -3283 289913 303275 290223
rect -3283 281213 303275 281523
rect -3283 279353 303275 279663
rect -3283 277493 303275 277803
rect -3283 275633 303275 275943
rect -3283 273773 303275 274083
rect -3283 271913 303275 272223
rect -3283 263213 303275 263523
rect -3283 261353 303275 261663
rect -3283 259493 303275 259803
rect -3283 257633 303275 257943
rect -3283 255773 303275 256083
rect -3283 253913 303275 254223
rect -3283 245213 303275 245523
rect -3283 243353 303275 243663
rect -3283 241493 303275 241803
rect -3283 239633 303275 239943
rect -3283 237773 303275 238083
rect -3283 235913 303275 236223
rect -3283 227213 303275 227523
rect -3283 225353 303275 225663
rect -3283 223493 303275 223803
rect -3283 221633 303275 221943
rect -3283 219773 303275 220083
rect -3283 217913 303275 218223
rect -3283 209213 303275 209523
rect -3283 207353 303275 207663
rect -3283 205493 303275 205803
rect -3283 203633 303275 203943
rect -3283 201773 303275 202083
rect -3283 199913 303275 200223
rect -3283 191213 303275 191523
rect -3283 189353 303275 189663
rect -3283 187493 303275 187803
rect -3283 185633 303275 185943
rect -3283 183773 303275 184083
rect -3283 181913 303275 182223
rect -3283 173213 303275 173523
rect -3283 171353 303275 171663
rect -3283 169493 303275 169803
rect -3283 167633 303275 167943
rect -3283 165773 303275 166083
rect -3283 163913 303275 164223
rect -3283 155213 303275 155523
rect -3283 153353 303275 153663
rect -3283 151493 303275 151803
rect -3283 149633 303275 149943
rect -3283 147773 303275 148083
rect -3283 145913 303275 146223
rect -3283 137213 303275 137523
rect -3283 135353 303275 135663
rect -3283 133493 303275 133803
rect -3283 131633 303275 131943
rect -3283 129773 303275 130083
rect -3283 127913 303275 128223
rect -3283 119213 303275 119523
rect -3283 117353 303275 117663
rect -3283 115493 303275 115803
rect -3283 113633 303275 113943
rect -3283 111773 303275 112083
rect -3283 109913 303275 110223
rect -3283 101213 303275 101523
rect -3283 99353 303275 99663
rect -3283 97493 303275 97803
rect -3283 95633 303275 95943
rect -3283 93773 303275 94083
rect -3283 91913 303275 92223
rect -3283 83213 303275 83523
rect -3283 81353 303275 81663
rect -3283 79493 303275 79803
rect -3283 77633 303275 77943
rect -3283 75773 303275 76083
rect -3283 73913 303275 74223
rect -3283 65213 303275 65523
rect -3283 63353 303275 63663
rect -3283 61493 303275 61803
rect -3283 59633 303275 59943
rect -3283 57773 303275 58083
rect -3283 55913 303275 56223
rect -3283 47213 303275 47523
rect -3283 45353 303275 45663
rect -3283 43493 303275 43803
rect -3283 41633 303275 41943
rect -3283 39773 303275 40083
rect -3283 37913 303275 38223
rect -3283 29213 303275 29523
rect -3283 27353 303275 27663
rect -3283 25493 303275 25803
rect -3283 23633 303275 23943
rect -3283 21773 303275 22083
rect -3283 19913 303275 20223
rect -3283 11213 303275 11523
rect -3283 9353 303275 9663
rect -3283 7493 303275 7803
rect -3283 5633 303275 5943
rect -3283 3773 303275 4083
rect -3283 1913 303275 2223
rect -883 13 300875 323
rect -1363 -467 301355 -157
rect -1843 -947 301835 -637
rect -2323 -1427 302315 -1117
rect -2803 -1907 302795 -1597
rect -3283 -2387 303275 -2077
<< labels >>
rlabel metal3 s 299760 2884 300480 2996 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 299760 195188 300480 195300 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 299760 217812 300480 217924 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 299760 240436 300480 240548 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 299760 263060 300480 263172 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 299760 285684 300480 285796 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 286692 299760 286804 300480 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 253540 299760 253652 300480 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 220388 299760 220500 300480 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 187236 299760 187348 300480 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 154084 299760 154196 300480 6 io_in[19]
port 11 nsew signal input
rlabel metal3 s 299760 19852 300480 19964 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 120932 299760 121044 300480 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 87780 299760 87892 300480 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 54628 299760 54740 300480 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 21476 299760 21588 300480 6 io_in[23]
port 16 nsew signal input
rlabel metal3 s -480 291284 240 291396 4 io_in[24]
port 17 nsew signal input
rlabel metal3 s -480 269108 240 269220 4 io_in[25]
port 18 nsew signal input
rlabel metal3 s -480 246932 240 247044 4 io_in[26]
port 19 nsew signal input
rlabel metal3 s -480 224756 240 224868 4 io_in[27]
port 20 nsew signal input
rlabel metal3 s -480 202580 240 202692 4 io_in[28]
port 21 nsew signal input
rlabel metal3 s -480 180404 240 180516 4 io_in[29]
port 22 nsew signal input
rlabel metal3 s 299760 36820 300480 36932 6 io_in[2]
port 23 nsew signal input
rlabel metal3 s -480 158228 240 158340 4 io_in[30]
port 24 nsew signal input
rlabel metal3 s -480 136052 240 136164 4 io_in[31]
port 25 nsew signal input
rlabel metal3 s -480 113876 240 113988 4 io_in[32]
port 26 nsew signal input
rlabel metal3 s -480 91700 240 91812 4 io_in[33]
port 27 nsew signal input
rlabel metal3 s -480 69524 240 69636 4 io_in[34]
port 28 nsew signal input
rlabel metal3 s -480 47348 240 47460 4 io_in[35]
port 29 nsew signal input
rlabel metal3 s -480 30716 240 30828 4 io_in[36]
port 30 nsew signal input
rlabel metal3 s -480 14084 240 14196 4 io_in[37]
port 31 nsew signal input
rlabel metal3 s 299760 53788 300480 53900 6 io_in[3]
port 32 nsew signal input
rlabel metal3 s 299760 70756 300480 70868 6 io_in[4]
port 33 nsew signal input
rlabel metal3 s 299760 87724 300480 87836 6 io_in[5]
port 34 nsew signal input
rlabel metal3 s 299760 104692 300480 104804 6 io_in[6]
port 35 nsew signal input
rlabel metal3 s 299760 127316 300480 127428 6 io_in[7]
port 36 nsew signal input
rlabel metal3 s 299760 149940 300480 150052 6 io_in[8]
port 37 nsew signal input
rlabel metal3 s 299760 172564 300480 172676 6 io_in[9]
port 38 nsew signal input
rlabel metal3 s 299760 14196 300480 14308 6 io_oeb[0]
port 39 nsew signal output
rlabel metal3 s 299760 206500 300480 206612 6 io_oeb[10]
port 40 nsew signal output
rlabel metal3 s 299760 229124 300480 229236 6 io_oeb[11]
port 41 nsew signal output
rlabel metal3 s 299760 251748 300480 251860 6 io_oeb[12]
port 42 nsew signal output
rlabel metal3 s 299760 274372 300480 274484 6 io_oeb[13]
port 43 nsew signal output
rlabel metal3 s 299760 296996 300480 297108 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 270116 299760 270228 300480 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 236964 299760 237076 300480 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 203812 299760 203924 300480 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 170660 299760 170772 300480 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 137508 299760 137620 300480 6 io_oeb[19]
port 49 nsew signal output
rlabel metal3 s 299760 31164 300480 31276 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 104356 299760 104468 300480 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 71204 299760 71316 300480 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 38052 299760 38164 300480 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 4900 299760 5012 300480 6 io_oeb[23]
port 54 nsew signal output
rlabel metal3 s -480 280196 240 280308 4 io_oeb[24]
port 55 nsew signal output
rlabel metal3 s -480 258020 240 258132 4 io_oeb[25]
port 56 nsew signal output
rlabel metal3 s -480 235844 240 235956 4 io_oeb[26]
port 57 nsew signal output
rlabel metal3 s -480 213668 240 213780 4 io_oeb[27]
port 58 nsew signal output
rlabel metal3 s -480 191492 240 191604 4 io_oeb[28]
port 59 nsew signal output
rlabel metal3 s -480 169316 240 169428 4 io_oeb[29]
port 60 nsew signal output
rlabel metal3 s 299760 48132 300480 48244 6 io_oeb[2]
port 61 nsew signal output
rlabel metal3 s -480 147140 240 147252 4 io_oeb[30]
port 62 nsew signal output
rlabel metal3 s -480 124964 240 125076 4 io_oeb[31]
port 63 nsew signal output
rlabel metal3 s -480 102788 240 102900 4 io_oeb[32]
port 64 nsew signal output
rlabel metal3 s -480 80612 240 80724 4 io_oeb[33]
port 65 nsew signal output
rlabel metal3 s -480 58436 240 58548 4 io_oeb[34]
port 66 nsew signal output
rlabel metal3 s -480 36260 240 36372 4 io_oeb[35]
port 67 nsew signal output
rlabel metal3 s -480 19628 240 19740 4 io_oeb[36]
port 68 nsew signal output
rlabel metal3 s -480 2996 240 3108 4 io_oeb[37]
port 69 nsew signal output
rlabel metal3 s 299760 65100 300480 65212 6 io_oeb[3]
port 70 nsew signal output
rlabel metal3 s 299760 82068 300480 82180 6 io_oeb[4]
port 71 nsew signal output
rlabel metal3 s 299760 99036 300480 99148 6 io_oeb[5]
port 72 nsew signal output
rlabel metal3 s 299760 116004 300480 116116 6 io_oeb[6]
port 73 nsew signal output
rlabel metal3 s 299760 138628 300480 138740 6 io_oeb[7]
port 74 nsew signal output
rlabel metal3 s 299760 161252 300480 161364 6 io_oeb[8]
port 75 nsew signal output
rlabel metal3 s 299760 183876 300480 183988 6 io_oeb[9]
port 76 nsew signal output
rlabel metal3 s 299760 8540 300480 8652 6 io_out[0]
port 77 nsew signal output
rlabel metal3 s 299760 200844 300480 200956 6 io_out[10]
port 78 nsew signal output
rlabel metal3 s 299760 223468 300480 223580 6 io_out[11]
port 79 nsew signal output
rlabel metal3 s 299760 246092 300480 246204 6 io_out[12]
port 80 nsew signal output
rlabel metal3 s 299760 268716 300480 268828 6 io_out[13]
port 81 nsew signal output
rlabel metal3 s 299760 291340 300480 291452 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 278404 299760 278516 300480 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 245252 299760 245364 300480 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 212100 299760 212212 300480 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 178948 299760 179060 300480 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 145796 299760 145908 300480 6 io_out[19]
port 87 nsew signal output
rlabel metal3 s 299760 25508 300480 25620 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 112644 299760 112756 300480 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 79492 299760 79604 300480 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 46340 299760 46452 300480 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 13188 299760 13300 300480 6 io_out[23]
port 92 nsew signal output
rlabel metal3 s -480 285740 240 285852 4 io_out[24]
port 93 nsew signal output
rlabel metal3 s -480 263564 240 263676 4 io_out[25]
port 94 nsew signal output
rlabel metal3 s -480 241388 240 241500 4 io_out[26]
port 95 nsew signal output
rlabel metal3 s -480 219212 240 219324 4 io_out[27]
port 96 nsew signal output
rlabel metal3 s -480 197036 240 197148 4 io_out[28]
port 97 nsew signal output
rlabel metal3 s -480 174860 240 174972 4 io_out[29]
port 98 nsew signal output
rlabel metal3 s 299760 42476 300480 42588 6 io_out[2]
port 99 nsew signal output
rlabel metal3 s -480 152684 240 152796 4 io_out[30]
port 100 nsew signal output
rlabel metal3 s -480 130508 240 130620 4 io_out[31]
port 101 nsew signal output
rlabel metal3 s -480 108332 240 108444 4 io_out[32]
port 102 nsew signal output
rlabel metal3 s -480 86156 240 86268 4 io_out[33]
port 103 nsew signal output
rlabel metal3 s -480 63980 240 64092 4 io_out[34]
port 104 nsew signal output
rlabel metal3 s -480 41804 240 41916 4 io_out[35]
port 105 nsew signal output
rlabel metal3 s -480 25172 240 25284 4 io_out[36]
port 106 nsew signal output
rlabel metal3 s -480 8540 240 8652 4 io_out[37]
port 107 nsew signal output
rlabel metal3 s 299760 59444 300480 59556 6 io_out[3]
port 108 nsew signal output
rlabel metal3 s 299760 76412 300480 76524 6 io_out[4]
port 109 nsew signal output
rlabel metal3 s 299760 93380 300480 93492 6 io_out[5]
port 110 nsew signal output
rlabel metal3 s 299760 110348 300480 110460 6 io_out[6]
port 111 nsew signal output
rlabel metal3 s 299760 132972 300480 133084 6 io_out[7]
port 112 nsew signal output
rlabel metal3 s 299760 155596 300480 155708 6 io_out[8]
port 113 nsew signal output
rlabel metal3 s 299760 178220 300480 178332 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 71260 -480 71372 240 8 la_data_in[0]
port 115 nsew signal input
rlabel metal2 s 88060 -480 88172 240 8 la_data_in[10]
port 116 nsew signal input
rlabel metal2 s 89740 -480 89852 240 8 la_data_in[11]
port 117 nsew signal input
rlabel metal2 s 91420 -480 91532 240 8 la_data_in[12]
port 118 nsew signal input
rlabel metal2 s 93100 -480 93212 240 8 la_data_in[13]
port 119 nsew signal input
rlabel metal2 s 94780 -480 94892 240 8 la_data_in[14]
port 120 nsew signal input
rlabel metal2 s 96460 -480 96572 240 8 la_data_in[15]
port 121 nsew signal input
rlabel metal2 s 98140 -480 98252 240 8 la_data_in[16]
port 122 nsew signal input
rlabel metal2 s 99820 -480 99932 240 8 la_data_in[17]
port 123 nsew signal input
rlabel metal2 s 101500 -480 101612 240 8 la_data_in[18]
port 124 nsew signal input
rlabel metal2 s 103180 -480 103292 240 8 la_data_in[19]
port 125 nsew signal input
rlabel metal2 s 72940 -480 73052 240 8 la_data_in[1]
port 126 nsew signal input
rlabel metal2 s 104860 -480 104972 240 8 la_data_in[20]
port 127 nsew signal input
rlabel metal2 s 106540 -480 106652 240 8 la_data_in[21]
port 128 nsew signal input
rlabel metal2 s 108220 -480 108332 240 8 la_data_in[22]
port 129 nsew signal input
rlabel metal2 s 109900 -480 110012 240 8 la_data_in[23]
port 130 nsew signal input
rlabel metal2 s 111580 -480 111692 240 8 la_data_in[24]
port 131 nsew signal input
rlabel metal2 s 113260 -480 113372 240 8 la_data_in[25]
port 132 nsew signal input
rlabel metal2 s 114940 -480 115052 240 8 la_data_in[26]
port 133 nsew signal input
rlabel metal2 s 116620 -480 116732 240 8 la_data_in[27]
port 134 nsew signal input
rlabel metal2 s 118300 -480 118412 240 8 la_data_in[28]
port 135 nsew signal input
rlabel metal2 s 119980 -480 120092 240 8 la_data_in[29]
port 136 nsew signal input
rlabel metal2 s 74620 -480 74732 240 8 la_data_in[2]
port 137 nsew signal input
rlabel metal2 s 121660 -480 121772 240 8 la_data_in[30]
port 138 nsew signal input
rlabel metal2 s 123340 -480 123452 240 8 la_data_in[31]
port 139 nsew signal input
rlabel metal2 s 125020 -480 125132 240 8 la_data_in[32]
port 140 nsew signal input
rlabel metal2 s 126700 -480 126812 240 8 la_data_in[33]
port 141 nsew signal input
rlabel metal2 s 128380 -480 128492 240 8 la_data_in[34]
port 142 nsew signal input
rlabel metal2 s 130060 -480 130172 240 8 la_data_in[35]
port 143 nsew signal input
rlabel metal2 s 131740 -480 131852 240 8 la_data_in[36]
port 144 nsew signal input
rlabel metal2 s 133420 -480 133532 240 8 la_data_in[37]
port 145 nsew signal input
rlabel metal2 s 135100 -480 135212 240 8 la_data_in[38]
port 146 nsew signal input
rlabel metal2 s 136780 -480 136892 240 8 la_data_in[39]
port 147 nsew signal input
rlabel metal2 s 76300 -480 76412 240 8 la_data_in[3]
port 148 nsew signal input
rlabel metal2 s 138460 -480 138572 240 8 la_data_in[40]
port 149 nsew signal input
rlabel metal2 s 140140 -480 140252 240 8 la_data_in[41]
port 150 nsew signal input
rlabel metal2 s 141820 -480 141932 240 8 la_data_in[42]
port 151 nsew signal input
rlabel metal2 s 143500 -480 143612 240 8 la_data_in[43]
port 152 nsew signal input
rlabel metal2 s 145180 -480 145292 240 8 la_data_in[44]
port 153 nsew signal input
rlabel metal2 s 146860 -480 146972 240 8 la_data_in[45]
port 154 nsew signal input
rlabel metal2 s 148540 -480 148652 240 8 la_data_in[46]
port 155 nsew signal input
rlabel metal2 s 150220 -480 150332 240 8 la_data_in[47]
port 156 nsew signal input
rlabel metal2 s 151900 -480 152012 240 8 la_data_in[48]
port 157 nsew signal input
rlabel metal2 s 153580 -480 153692 240 8 la_data_in[49]
port 158 nsew signal input
rlabel metal2 s 77980 -480 78092 240 8 la_data_in[4]
port 159 nsew signal input
rlabel metal2 s 155260 -480 155372 240 8 la_data_in[50]
port 160 nsew signal input
rlabel metal2 s 156940 -480 157052 240 8 la_data_in[51]
port 161 nsew signal input
rlabel metal2 s 158620 -480 158732 240 8 la_data_in[52]
port 162 nsew signal input
rlabel metal2 s 160300 -480 160412 240 8 la_data_in[53]
port 163 nsew signal input
rlabel metal2 s 161980 -480 162092 240 8 la_data_in[54]
port 164 nsew signal input
rlabel metal2 s 163660 -480 163772 240 8 la_data_in[55]
port 165 nsew signal input
rlabel metal2 s 165340 -480 165452 240 8 la_data_in[56]
port 166 nsew signal input
rlabel metal2 s 167020 -480 167132 240 8 la_data_in[57]
port 167 nsew signal input
rlabel metal2 s 168700 -480 168812 240 8 la_data_in[58]
port 168 nsew signal input
rlabel metal2 s 170380 -480 170492 240 8 la_data_in[59]
port 169 nsew signal input
rlabel metal2 s 79660 -480 79772 240 8 la_data_in[5]
port 170 nsew signal input
rlabel metal2 s 172060 -480 172172 240 8 la_data_in[60]
port 171 nsew signal input
rlabel metal2 s 173740 -480 173852 240 8 la_data_in[61]
port 172 nsew signal input
rlabel metal2 s 175420 -480 175532 240 8 la_data_in[62]
port 173 nsew signal input
rlabel metal2 s 177100 -480 177212 240 8 la_data_in[63]
port 174 nsew signal input
rlabel metal2 s 81340 -480 81452 240 8 la_data_in[6]
port 175 nsew signal input
rlabel metal2 s 83020 -480 83132 240 8 la_data_in[7]
port 176 nsew signal input
rlabel metal2 s 84700 -480 84812 240 8 la_data_in[8]
port 177 nsew signal input
rlabel metal2 s 86380 -480 86492 240 8 la_data_in[9]
port 178 nsew signal input
rlabel metal2 s 71820 -480 71932 240 8 la_data_out[0]
port 179 nsew signal output
rlabel metal2 s 88620 -480 88732 240 8 la_data_out[10]
port 180 nsew signal output
rlabel metal2 s 90300 -480 90412 240 8 la_data_out[11]
port 181 nsew signal output
rlabel metal2 s 91980 -480 92092 240 8 la_data_out[12]
port 182 nsew signal output
rlabel metal2 s 93660 -480 93772 240 8 la_data_out[13]
port 183 nsew signal output
rlabel metal2 s 95340 -480 95452 240 8 la_data_out[14]
port 184 nsew signal output
rlabel metal2 s 97020 -480 97132 240 8 la_data_out[15]
port 185 nsew signal output
rlabel metal2 s 98700 -480 98812 240 8 la_data_out[16]
port 186 nsew signal output
rlabel metal2 s 100380 -480 100492 240 8 la_data_out[17]
port 187 nsew signal output
rlabel metal2 s 102060 -480 102172 240 8 la_data_out[18]
port 188 nsew signal output
rlabel metal2 s 103740 -480 103852 240 8 la_data_out[19]
port 189 nsew signal output
rlabel metal2 s 73500 -480 73612 240 8 la_data_out[1]
port 190 nsew signal output
rlabel metal2 s 105420 -480 105532 240 8 la_data_out[20]
port 191 nsew signal output
rlabel metal2 s 107100 -480 107212 240 8 la_data_out[21]
port 192 nsew signal output
rlabel metal2 s 108780 -480 108892 240 8 la_data_out[22]
port 193 nsew signal output
rlabel metal2 s 110460 -480 110572 240 8 la_data_out[23]
port 194 nsew signal output
rlabel metal2 s 112140 -480 112252 240 8 la_data_out[24]
port 195 nsew signal output
rlabel metal2 s 113820 -480 113932 240 8 la_data_out[25]
port 196 nsew signal output
rlabel metal2 s 115500 -480 115612 240 8 la_data_out[26]
port 197 nsew signal output
rlabel metal2 s 117180 -480 117292 240 8 la_data_out[27]
port 198 nsew signal output
rlabel metal2 s 118860 -480 118972 240 8 la_data_out[28]
port 199 nsew signal output
rlabel metal2 s 120540 -480 120652 240 8 la_data_out[29]
port 200 nsew signal output
rlabel metal2 s 75180 -480 75292 240 8 la_data_out[2]
port 201 nsew signal output
rlabel metal2 s 122220 -480 122332 240 8 la_data_out[30]
port 202 nsew signal output
rlabel metal2 s 123900 -480 124012 240 8 la_data_out[31]
port 203 nsew signal output
rlabel metal2 s 125580 -480 125692 240 8 la_data_out[32]
port 204 nsew signal output
rlabel metal2 s 127260 -480 127372 240 8 la_data_out[33]
port 205 nsew signal output
rlabel metal2 s 128940 -480 129052 240 8 la_data_out[34]
port 206 nsew signal output
rlabel metal2 s 130620 -480 130732 240 8 la_data_out[35]
port 207 nsew signal output
rlabel metal2 s 132300 -480 132412 240 8 la_data_out[36]
port 208 nsew signal output
rlabel metal2 s 133980 -480 134092 240 8 la_data_out[37]
port 209 nsew signal output
rlabel metal2 s 135660 -480 135772 240 8 la_data_out[38]
port 210 nsew signal output
rlabel metal2 s 137340 -480 137452 240 8 la_data_out[39]
port 211 nsew signal output
rlabel metal2 s 76860 -480 76972 240 8 la_data_out[3]
port 212 nsew signal output
rlabel metal2 s 139020 -480 139132 240 8 la_data_out[40]
port 213 nsew signal output
rlabel metal2 s 140700 -480 140812 240 8 la_data_out[41]
port 214 nsew signal output
rlabel metal2 s 142380 -480 142492 240 8 la_data_out[42]
port 215 nsew signal output
rlabel metal2 s 144060 -480 144172 240 8 la_data_out[43]
port 216 nsew signal output
rlabel metal2 s 145740 -480 145852 240 8 la_data_out[44]
port 217 nsew signal output
rlabel metal2 s 147420 -480 147532 240 8 la_data_out[45]
port 218 nsew signal output
rlabel metal2 s 149100 -480 149212 240 8 la_data_out[46]
port 219 nsew signal output
rlabel metal2 s 150780 -480 150892 240 8 la_data_out[47]
port 220 nsew signal output
rlabel metal2 s 152460 -480 152572 240 8 la_data_out[48]
port 221 nsew signal output
rlabel metal2 s 154140 -480 154252 240 8 la_data_out[49]
port 222 nsew signal output
rlabel metal2 s 78540 -480 78652 240 8 la_data_out[4]
port 223 nsew signal output
rlabel metal2 s 155820 -480 155932 240 8 la_data_out[50]
port 224 nsew signal output
rlabel metal2 s 157500 -480 157612 240 8 la_data_out[51]
port 225 nsew signal output
rlabel metal2 s 159180 -480 159292 240 8 la_data_out[52]
port 226 nsew signal output
rlabel metal2 s 160860 -480 160972 240 8 la_data_out[53]
port 227 nsew signal output
rlabel metal2 s 162540 -480 162652 240 8 la_data_out[54]
port 228 nsew signal output
rlabel metal2 s 164220 -480 164332 240 8 la_data_out[55]
port 229 nsew signal output
rlabel metal2 s 165900 -480 166012 240 8 la_data_out[56]
port 230 nsew signal output
rlabel metal2 s 167580 -480 167692 240 8 la_data_out[57]
port 231 nsew signal output
rlabel metal2 s 169260 -480 169372 240 8 la_data_out[58]
port 232 nsew signal output
rlabel metal2 s 170940 -480 171052 240 8 la_data_out[59]
port 233 nsew signal output
rlabel metal2 s 80220 -480 80332 240 8 la_data_out[5]
port 234 nsew signal output
rlabel metal2 s 172620 -480 172732 240 8 la_data_out[60]
port 235 nsew signal output
rlabel metal2 s 174300 -480 174412 240 8 la_data_out[61]
port 236 nsew signal output
rlabel metal2 s 175980 -480 176092 240 8 la_data_out[62]
port 237 nsew signal output
rlabel metal2 s 177660 -480 177772 240 8 la_data_out[63]
port 238 nsew signal output
rlabel metal2 s 81900 -480 82012 240 8 la_data_out[6]
port 239 nsew signal output
rlabel metal2 s 83580 -480 83692 240 8 la_data_out[7]
port 240 nsew signal output
rlabel metal2 s 85260 -480 85372 240 8 la_data_out[8]
port 241 nsew signal output
rlabel metal2 s 86940 -480 87052 240 8 la_data_out[9]
port 242 nsew signal output
rlabel metal2 s 72380 -480 72492 240 8 la_oenb[0]
port 243 nsew signal input
rlabel metal2 s 89180 -480 89292 240 8 la_oenb[10]
port 244 nsew signal input
rlabel metal2 s 90860 -480 90972 240 8 la_oenb[11]
port 245 nsew signal input
rlabel metal2 s 92540 -480 92652 240 8 la_oenb[12]
port 246 nsew signal input
rlabel metal2 s 94220 -480 94332 240 8 la_oenb[13]
port 247 nsew signal input
rlabel metal2 s 95900 -480 96012 240 8 la_oenb[14]
port 248 nsew signal input
rlabel metal2 s 97580 -480 97692 240 8 la_oenb[15]
port 249 nsew signal input
rlabel metal2 s 99260 -480 99372 240 8 la_oenb[16]
port 250 nsew signal input
rlabel metal2 s 100940 -480 101052 240 8 la_oenb[17]
port 251 nsew signal input
rlabel metal2 s 102620 -480 102732 240 8 la_oenb[18]
port 252 nsew signal input
rlabel metal2 s 104300 -480 104412 240 8 la_oenb[19]
port 253 nsew signal input
rlabel metal2 s 74060 -480 74172 240 8 la_oenb[1]
port 254 nsew signal input
rlabel metal2 s 105980 -480 106092 240 8 la_oenb[20]
port 255 nsew signal input
rlabel metal2 s 107660 -480 107772 240 8 la_oenb[21]
port 256 nsew signal input
rlabel metal2 s 109340 -480 109452 240 8 la_oenb[22]
port 257 nsew signal input
rlabel metal2 s 111020 -480 111132 240 8 la_oenb[23]
port 258 nsew signal input
rlabel metal2 s 112700 -480 112812 240 8 la_oenb[24]
port 259 nsew signal input
rlabel metal2 s 114380 -480 114492 240 8 la_oenb[25]
port 260 nsew signal input
rlabel metal2 s 116060 -480 116172 240 8 la_oenb[26]
port 261 nsew signal input
rlabel metal2 s 117740 -480 117852 240 8 la_oenb[27]
port 262 nsew signal input
rlabel metal2 s 119420 -480 119532 240 8 la_oenb[28]
port 263 nsew signal input
rlabel metal2 s 121100 -480 121212 240 8 la_oenb[29]
port 264 nsew signal input
rlabel metal2 s 75740 -480 75852 240 8 la_oenb[2]
port 265 nsew signal input
rlabel metal2 s 122780 -480 122892 240 8 la_oenb[30]
port 266 nsew signal input
rlabel metal2 s 124460 -480 124572 240 8 la_oenb[31]
port 267 nsew signal input
rlabel metal2 s 126140 -480 126252 240 8 la_oenb[32]
port 268 nsew signal input
rlabel metal2 s 127820 -480 127932 240 8 la_oenb[33]
port 269 nsew signal input
rlabel metal2 s 129500 -480 129612 240 8 la_oenb[34]
port 270 nsew signal input
rlabel metal2 s 131180 -480 131292 240 8 la_oenb[35]
port 271 nsew signal input
rlabel metal2 s 132860 -480 132972 240 8 la_oenb[36]
port 272 nsew signal input
rlabel metal2 s 134540 -480 134652 240 8 la_oenb[37]
port 273 nsew signal input
rlabel metal2 s 136220 -480 136332 240 8 la_oenb[38]
port 274 nsew signal input
rlabel metal2 s 137900 -480 138012 240 8 la_oenb[39]
port 275 nsew signal input
rlabel metal2 s 77420 -480 77532 240 8 la_oenb[3]
port 276 nsew signal input
rlabel metal2 s 139580 -480 139692 240 8 la_oenb[40]
port 277 nsew signal input
rlabel metal2 s 141260 -480 141372 240 8 la_oenb[41]
port 278 nsew signal input
rlabel metal2 s 142940 -480 143052 240 8 la_oenb[42]
port 279 nsew signal input
rlabel metal2 s 144620 -480 144732 240 8 la_oenb[43]
port 280 nsew signal input
rlabel metal2 s 146300 -480 146412 240 8 la_oenb[44]
port 281 nsew signal input
rlabel metal2 s 147980 -480 148092 240 8 la_oenb[45]
port 282 nsew signal input
rlabel metal2 s 149660 -480 149772 240 8 la_oenb[46]
port 283 nsew signal input
rlabel metal2 s 151340 -480 151452 240 8 la_oenb[47]
port 284 nsew signal input
rlabel metal2 s 153020 -480 153132 240 8 la_oenb[48]
port 285 nsew signal input
rlabel metal2 s 154700 -480 154812 240 8 la_oenb[49]
port 286 nsew signal input
rlabel metal2 s 79100 -480 79212 240 8 la_oenb[4]
port 287 nsew signal input
rlabel metal2 s 156380 -480 156492 240 8 la_oenb[50]
port 288 nsew signal input
rlabel metal2 s 158060 -480 158172 240 8 la_oenb[51]
port 289 nsew signal input
rlabel metal2 s 159740 -480 159852 240 8 la_oenb[52]
port 290 nsew signal input
rlabel metal2 s 161420 -480 161532 240 8 la_oenb[53]
port 291 nsew signal input
rlabel metal2 s 163100 -480 163212 240 8 la_oenb[54]
port 292 nsew signal input
rlabel metal2 s 164780 -480 164892 240 8 la_oenb[55]
port 293 nsew signal input
rlabel metal2 s 166460 -480 166572 240 8 la_oenb[56]
port 294 nsew signal input
rlabel metal2 s 168140 -480 168252 240 8 la_oenb[57]
port 295 nsew signal input
rlabel metal2 s 169820 -480 169932 240 8 la_oenb[58]
port 296 nsew signal input
rlabel metal2 s 171500 -480 171612 240 8 la_oenb[59]
port 297 nsew signal input
rlabel metal2 s 80780 -480 80892 240 8 la_oenb[5]
port 298 nsew signal input
rlabel metal2 s 173180 -480 173292 240 8 la_oenb[60]
port 299 nsew signal input
rlabel metal2 s 174860 -480 174972 240 8 la_oenb[61]
port 300 nsew signal input
rlabel metal2 s 176540 -480 176652 240 8 la_oenb[62]
port 301 nsew signal input
rlabel metal2 s 178220 -480 178332 240 8 la_oenb[63]
port 302 nsew signal input
rlabel metal2 s 82460 -480 82572 240 8 la_oenb[6]
port 303 nsew signal input
rlabel metal2 s 84140 -480 84252 240 8 la_oenb[7]
port 304 nsew signal input
rlabel metal2 s 85820 -480 85932 240 8 la_oenb[8]
port 305 nsew signal input
rlabel metal2 s 87500 -480 87612 240 8 la_oenb[9]
port 306 nsew signal input
rlabel metal2 s 286300 -480 286412 240 8 user_clock2
port 307 nsew signal input
rlabel metal2 s 286860 -480 286972 240 8 user_irq[0]
port 308 nsew signal output
rlabel metal2 s 287420 -480 287532 240 8 user_irq[1]
port 309 nsew signal output
rlabel metal2 s 287980 -480 288092 240 8 user_irq[2]
port 310 nsew signal output
rlabel metal4 s -883 13 -573 299867 4 vccd1
port 311 nsew power bidirectional
rlabel metal5 s -883 13 300875 323 6 vccd1
port 311 nsew power bidirectional
rlabel metal5 s -883 299557 300875 299867 6 vccd1
port 311 nsew power bidirectional
rlabel metal4 s 300565 13 300875 299867 6 vccd1
port 311 nsew power bidirectional
rlabel metal4 s 1017 -2387 1327 302267 6 vccd1
port 311 nsew power bidirectional
rlabel metal4 s 19017 -2387 19327 302267 6 vccd1
port 311 nsew power bidirectional
rlabel metal4 s 37017 -2387 37327 82289 6 vccd1
port 311 nsew power bidirectional
rlabel metal4 s 37017 94967 37327 302267 6 vccd1
port 311 nsew power bidirectional
rlabel metal4 s 55017 -2387 55327 51721 6 vccd1
port 311 nsew power bidirectional
rlabel metal4 s 55017 59415 55327 302267 6 vccd1
port 311 nsew power bidirectional
rlabel metal4 s 73017 -2387 73327 302267 6 vccd1
port 311 nsew power bidirectional
rlabel metal4 s 91017 -2387 91327 302267 6 vccd1
port 311 nsew power bidirectional
rlabel metal4 s 109017 -2387 109327 302267 6 vccd1
port 311 nsew power bidirectional
rlabel metal4 s 127017 -2387 127327 302267 6 vccd1
port 311 nsew power bidirectional
rlabel metal4 s 145017 -2387 145327 302267 6 vccd1
port 311 nsew power bidirectional
rlabel metal4 s 163017 -2387 163327 302267 6 vccd1
port 311 nsew power bidirectional
rlabel metal4 s 181017 -2387 181327 302267 6 vccd1
port 311 nsew power bidirectional
rlabel metal4 s 199017 -2387 199327 302267 6 vccd1
port 311 nsew power bidirectional
rlabel metal4 s 217017 -2387 217327 302267 6 vccd1
port 311 nsew power bidirectional
rlabel metal4 s 235017 -2387 235327 302267 6 vccd1
port 311 nsew power bidirectional
rlabel metal4 s 253017 -2387 253327 302267 6 vccd1
port 311 nsew power bidirectional
rlabel metal4 s 271017 -2387 271327 302267 6 vccd1
port 311 nsew power bidirectional
rlabel metal4 s 289017 -2387 289327 302267 6 vccd1
port 311 nsew power bidirectional
rlabel metal5 s -3283 1913 303275 2223 6 vccd1
port 311 nsew power bidirectional
rlabel metal5 s -3283 19913 303275 20223 6 vccd1
port 311 nsew power bidirectional
rlabel metal5 s -3283 37913 303275 38223 6 vccd1
port 311 nsew power bidirectional
rlabel metal5 s -3283 55913 303275 56223 6 vccd1
port 311 nsew power bidirectional
rlabel metal5 s -3283 73913 303275 74223 6 vccd1
port 311 nsew power bidirectional
rlabel metal5 s -3283 91913 303275 92223 6 vccd1
port 311 nsew power bidirectional
rlabel metal5 s -3283 109913 303275 110223 6 vccd1
port 311 nsew power bidirectional
rlabel metal5 s -3283 127913 303275 128223 6 vccd1
port 311 nsew power bidirectional
rlabel metal5 s -3283 145913 303275 146223 6 vccd1
port 311 nsew power bidirectional
rlabel metal5 s -3283 163913 303275 164223 6 vccd1
port 311 nsew power bidirectional
rlabel metal5 s -3283 181913 303275 182223 6 vccd1
port 311 nsew power bidirectional
rlabel metal5 s -3283 199913 303275 200223 6 vccd1
port 311 nsew power bidirectional
rlabel metal5 s -3283 217913 303275 218223 6 vccd1
port 311 nsew power bidirectional
rlabel metal5 s -3283 235913 303275 236223 6 vccd1
port 311 nsew power bidirectional
rlabel metal5 s -3283 253913 303275 254223 6 vccd1
port 311 nsew power bidirectional
rlabel metal5 s -3283 271913 303275 272223 6 vccd1
port 311 nsew power bidirectional
rlabel metal5 s -3283 289913 303275 290223 6 vccd1
port 311 nsew power bidirectional
rlabel metal4 s -1843 -947 -1533 300827 4 vccd2
port 312 nsew power bidirectional
rlabel metal5 s -1843 -947 301835 -637 8 vccd2
port 312 nsew power bidirectional
rlabel metal5 s -1843 300517 301835 300827 6 vccd2
port 312 nsew power bidirectional
rlabel metal4 s 301525 -947 301835 300827 6 vccd2
port 312 nsew power bidirectional
rlabel metal4 s 4737 -2387 5047 302267 6 vccd2
port 312 nsew power bidirectional
rlabel metal4 s 22737 -2387 23047 302267 6 vccd2
port 312 nsew power bidirectional
rlabel metal4 s 40737 -2387 41047 82289 6 vccd2
port 312 nsew power bidirectional
rlabel metal4 s 40737 94967 41047 302267 6 vccd2
port 312 nsew power bidirectional
rlabel metal4 s 58737 -2387 59047 51721 6 vccd2
port 312 nsew power bidirectional
rlabel metal4 s 58737 59415 59047 302267 6 vccd2
port 312 nsew power bidirectional
rlabel metal4 s 76737 -2387 77047 302267 6 vccd2
port 312 nsew power bidirectional
rlabel metal4 s 94737 -2387 95047 302267 6 vccd2
port 312 nsew power bidirectional
rlabel metal4 s 112737 -2387 113047 302267 6 vccd2
port 312 nsew power bidirectional
rlabel metal4 s 130737 -2387 131047 302267 6 vccd2
port 312 nsew power bidirectional
rlabel metal4 s 148737 -2387 149047 302267 6 vccd2
port 312 nsew power bidirectional
rlabel metal4 s 166737 -2387 167047 302267 6 vccd2
port 312 nsew power bidirectional
rlabel metal4 s 184737 -2387 185047 302267 6 vccd2
port 312 nsew power bidirectional
rlabel metal4 s 202737 -2387 203047 302267 6 vccd2
port 312 nsew power bidirectional
rlabel metal4 s 220737 -2387 221047 302267 6 vccd2
port 312 nsew power bidirectional
rlabel metal4 s 238737 -2387 239047 302267 6 vccd2
port 312 nsew power bidirectional
rlabel metal4 s 256737 -2387 257047 302267 6 vccd2
port 312 nsew power bidirectional
rlabel metal4 s 274737 -2387 275047 302267 6 vccd2
port 312 nsew power bidirectional
rlabel metal4 s 292737 -2387 293047 302267 6 vccd2
port 312 nsew power bidirectional
rlabel metal5 s -3283 5633 303275 5943 6 vccd2
port 312 nsew power bidirectional
rlabel metal5 s -3283 23633 303275 23943 6 vccd2
port 312 nsew power bidirectional
rlabel metal5 s -3283 41633 303275 41943 6 vccd2
port 312 nsew power bidirectional
rlabel metal5 s -3283 59633 303275 59943 6 vccd2
port 312 nsew power bidirectional
rlabel metal5 s -3283 77633 303275 77943 6 vccd2
port 312 nsew power bidirectional
rlabel metal5 s -3283 95633 303275 95943 6 vccd2
port 312 nsew power bidirectional
rlabel metal5 s -3283 113633 303275 113943 6 vccd2
port 312 nsew power bidirectional
rlabel metal5 s -3283 131633 303275 131943 6 vccd2
port 312 nsew power bidirectional
rlabel metal5 s -3283 149633 303275 149943 6 vccd2
port 312 nsew power bidirectional
rlabel metal5 s -3283 167633 303275 167943 6 vccd2
port 312 nsew power bidirectional
rlabel metal5 s -3283 185633 303275 185943 6 vccd2
port 312 nsew power bidirectional
rlabel metal5 s -3283 203633 303275 203943 6 vccd2
port 312 nsew power bidirectional
rlabel metal5 s -3283 221633 303275 221943 6 vccd2
port 312 nsew power bidirectional
rlabel metal5 s -3283 239633 303275 239943 6 vccd2
port 312 nsew power bidirectional
rlabel metal5 s -3283 257633 303275 257943 6 vccd2
port 312 nsew power bidirectional
rlabel metal5 s -3283 275633 303275 275943 6 vccd2
port 312 nsew power bidirectional
rlabel metal5 s -3283 293633 303275 293943 6 vccd2
port 312 nsew power bidirectional
rlabel metal4 s -2803 -1907 -2493 301787 4 vdda1
port 313 nsew power bidirectional
rlabel metal5 s -2803 -1907 302795 -1597 8 vdda1
port 313 nsew power bidirectional
rlabel metal5 s -2803 301477 302795 301787 6 vdda1
port 313 nsew power bidirectional
rlabel metal4 s 302485 -1907 302795 301787 6 vdda1
port 313 nsew power bidirectional
rlabel metal4 s 8457 -2387 8767 302267 6 vdda1
port 313 nsew power bidirectional
rlabel metal4 s 26457 -2387 26767 82289 6 vdda1
port 313 nsew power bidirectional
rlabel metal4 s 26457 94967 26767 302267 6 vdda1
port 313 nsew power bidirectional
rlabel metal4 s 44457 -2387 44767 51721 6 vdda1
port 313 nsew power bidirectional
rlabel metal4 s 44457 59415 44767 82289 6 vdda1
port 313 nsew power bidirectional
rlabel metal4 s 44457 94967 44767 302267 6 vdda1
port 313 nsew power bidirectional
rlabel metal4 s 62457 -2387 62767 302267 6 vdda1
port 313 nsew power bidirectional
rlabel metal4 s 80457 -2387 80767 302267 6 vdda1
port 313 nsew power bidirectional
rlabel metal4 s 98457 -2387 98767 302267 6 vdda1
port 313 nsew power bidirectional
rlabel metal4 s 116457 -2387 116767 302267 6 vdda1
port 313 nsew power bidirectional
rlabel metal4 s 134457 -2387 134767 302267 6 vdda1
port 313 nsew power bidirectional
rlabel metal4 s 152457 -2387 152767 302267 6 vdda1
port 313 nsew power bidirectional
rlabel metal4 s 170457 -2387 170767 302267 6 vdda1
port 313 nsew power bidirectional
rlabel metal4 s 188457 -2387 188767 302267 6 vdda1
port 313 nsew power bidirectional
rlabel metal4 s 206457 -2387 206767 302267 6 vdda1
port 313 nsew power bidirectional
rlabel metal4 s 224457 -2387 224767 302267 6 vdda1
port 313 nsew power bidirectional
rlabel metal4 s 242457 -2387 242767 302267 6 vdda1
port 313 nsew power bidirectional
rlabel metal4 s 260457 -2387 260767 302267 6 vdda1
port 313 nsew power bidirectional
rlabel metal4 s 278457 -2387 278767 302267 6 vdda1
port 313 nsew power bidirectional
rlabel metal4 s 296457 -2387 296767 302267 6 vdda1
port 313 nsew power bidirectional
rlabel metal5 s -3283 9353 303275 9663 6 vdda1
port 313 nsew power bidirectional
rlabel metal5 s -3283 27353 303275 27663 6 vdda1
port 313 nsew power bidirectional
rlabel metal5 s -3283 45353 303275 45663 6 vdda1
port 313 nsew power bidirectional
rlabel metal5 s -3283 63353 303275 63663 6 vdda1
port 313 nsew power bidirectional
rlabel metal5 s -3283 81353 303275 81663 6 vdda1
port 313 nsew power bidirectional
rlabel metal5 s -3283 99353 303275 99663 6 vdda1
port 313 nsew power bidirectional
rlabel metal5 s -3283 117353 303275 117663 6 vdda1
port 313 nsew power bidirectional
rlabel metal5 s -3283 135353 303275 135663 6 vdda1
port 313 nsew power bidirectional
rlabel metal5 s -3283 153353 303275 153663 6 vdda1
port 313 nsew power bidirectional
rlabel metal5 s -3283 171353 303275 171663 6 vdda1
port 313 nsew power bidirectional
rlabel metal5 s -3283 189353 303275 189663 6 vdda1
port 313 nsew power bidirectional
rlabel metal5 s -3283 207353 303275 207663 6 vdda1
port 313 nsew power bidirectional
rlabel metal5 s -3283 225353 303275 225663 6 vdda1
port 313 nsew power bidirectional
rlabel metal5 s -3283 243353 303275 243663 6 vdda1
port 313 nsew power bidirectional
rlabel metal5 s -3283 261353 303275 261663 6 vdda1
port 313 nsew power bidirectional
rlabel metal5 s -3283 279353 303275 279663 6 vdda1
port 313 nsew power bidirectional
rlabel metal5 s -3283 297353 303275 297663 6 vdda1
port 313 nsew power bidirectional
rlabel metal4 s -3283 -2387 -2973 302267 4 vssa1
port 314 nsew ground bidirectional
rlabel metal5 s -3283 -2387 303275 -2077 8 vssa1
port 314 nsew ground bidirectional
rlabel metal5 s -3283 301957 303275 302267 6 vssa1
port 314 nsew ground bidirectional
rlabel metal4 s 302965 -2387 303275 302267 6 vssa1
port 314 nsew ground bidirectional
rlabel metal4 s 10317 -2387 10627 302267 6 vssa1
port 314 nsew ground bidirectional
rlabel metal4 s 28317 -2387 28627 82289 6 vssa1
port 314 nsew ground bidirectional
rlabel metal4 s 28317 94967 28627 302267 6 vssa1
port 314 nsew ground bidirectional
rlabel metal4 s 46317 -2387 46627 51721 6 vssa1
port 314 nsew ground bidirectional
rlabel metal4 s 46317 59415 46627 302267 6 vssa1
port 314 nsew ground bidirectional
rlabel metal4 s 64317 -2387 64627 302267 6 vssa1
port 314 nsew ground bidirectional
rlabel metal4 s 82317 -2387 82627 302267 6 vssa1
port 314 nsew ground bidirectional
rlabel metal4 s 100317 -2387 100627 302267 6 vssa1
port 314 nsew ground bidirectional
rlabel metal4 s 118317 -2387 118627 302267 6 vssa1
port 314 nsew ground bidirectional
rlabel metal4 s 136317 -2387 136627 302267 6 vssa1
port 314 nsew ground bidirectional
rlabel metal4 s 154317 -2387 154627 302267 6 vssa1
port 314 nsew ground bidirectional
rlabel metal4 s 172317 -2387 172627 302267 6 vssa1
port 314 nsew ground bidirectional
rlabel metal4 s 190317 -2387 190627 302267 6 vssa1
port 314 nsew ground bidirectional
rlabel metal4 s 208317 -2387 208627 302267 6 vssa1
port 314 nsew ground bidirectional
rlabel metal4 s 226317 -2387 226627 302267 6 vssa1
port 314 nsew ground bidirectional
rlabel metal4 s 244317 -2387 244627 302267 6 vssa1
port 314 nsew ground bidirectional
rlabel metal4 s 262317 -2387 262627 302267 6 vssa1
port 314 nsew ground bidirectional
rlabel metal4 s 280317 -2387 280627 302267 6 vssa1
port 314 nsew ground bidirectional
rlabel metal4 s 298317 -2387 298627 302267 6 vssa1
port 314 nsew ground bidirectional
rlabel metal5 s -3283 11213 303275 11523 6 vssa1
port 314 nsew ground bidirectional
rlabel metal5 s -3283 29213 303275 29523 6 vssa1
port 314 nsew ground bidirectional
rlabel metal5 s -3283 47213 303275 47523 6 vssa1
port 314 nsew ground bidirectional
rlabel metal5 s -3283 65213 303275 65523 6 vssa1
port 314 nsew ground bidirectional
rlabel metal5 s -3283 83213 303275 83523 6 vssa1
port 314 nsew ground bidirectional
rlabel metal5 s -3283 101213 303275 101523 6 vssa1
port 314 nsew ground bidirectional
rlabel metal5 s -3283 119213 303275 119523 6 vssa1
port 314 nsew ground bidirectional
rlabel metal5 s -3283 137213 303275 137523 6 vssa1
port 314 nsew ground bidirectional
rlabel metal5 s -3283 155213 303275 155523 6 vssa1
port 314 nsew ground bidirectional
rlabel metal5 s -3283 173213 303275 173523 6 vssa1
port 314 nsew ground bidirectional
rlabel metal5 s -3283 191213 303275 191523 6 vssa1
port 314 nsew ground bidirectional
rlabel metal5 s -3283 209213 303275 209523 6 vssa1
port 314 nsew ground bidirectional
rlabel metal5 s -3283 227213 303275 227523 6 vssa1
port 314 nsew ground bidirectional
rlabel metal5 s -3283 245213 303275 245523 6 vssa1
port 314 nsew ground bidirectional
rlabel metal5 s -3283 263213 303275 263523 6 vssa1
port 314 nsew ground bidirectional
rlabel metal5 s -3283 281213 303275 281523 6 vssa1
port 314 nsew ground bidirectional
rlabel metal4 s -1363 -467 -1053 300347 4 vssd1
port 315 nsew ground bidirectional
rlabel metal5 s -1363 -467 301355 -157 8 vssd1
port 315 nsew ground bidirectional
rlabel metal5 s -1363 300037 301355 300347 6 vssd1
port 315 nsew ground bidirectional
rlabel metal4 s 301045 -467 301355 300347 6 vssd1
port 315 nsew ground bidirectional
rlabel metal4 s 2877 -2387 3187 302267 6 vssd1
port 315 nsew ground bidirectional
rlabel metal4 s 20877 -2387 21187 302267 6 vssd1
port 315 nsew ground bidirectional
rlabel metal4 s 38877 -2387 39187 82289 6 vssd1
port 315 nsew ground bidirectional
rlabel metal4 s 38877 94967 39187 302267 6 vssd1
port 315 nsew ground bidirectional
rlabel metal4 s 56877 -2387 57187 51721 6 vssd1
port 315 nsew ground bidirectional
rlabel metal4 s 56877 59415 57187 302267 6 vssd1
port 315 nsew ground bidirectional
rlabel metal4 s 74877 -2387 75187 302267 6 vssd1
port 315 nsew ground bidirectional
rlabel metal4 s 92877 -2387 93187 302267 6 vssd1
port 315 nsew ground bidirectional
rlabel metal4 s 110877 -2387 111187 302267 6 vssd1
port 315 nsew ground bidirectional
rlabel metal4 s 128877 -2387 129187 302267 6 vssd1
port 315 nsew ground bidirectional
rlabel metal4 s 146877 -2387 147187 302267 6 vssd1
port 315 nsew ground bidirectional
rlabel metal4 s 164877 -2387 165187 302267 6 vssd1
port 315 nsew ground bidirectional
rlabel metal4 s 182877 -2387 183187 302267 6 vssd1
port 315 nsew ground bidirectional
rlabel metal4 s 200877 -2387 201187 302267 6 vssd1
port 315 nsew ground bidirectional
rlabel metal4 s 218877 -2387 219187 302267 6 vssd1
port 315 nsew ground bidirectional
rlabel metal4 s 236877 -2387 237187 302267 6 vssd1
port 315 nsew ground bidirectional
rlabel metal4 s 254877 -2387 255187 302267 6 vssd1
port 315 nsew ground bidirectional
rlabel metal4 s 272877 -2387 273187 302267 6 vssd1
port 315 nsew ground bidirectional
rlabel metal4 s 290877 -2387 291187 302267 6 vssd1
port 315 nsew ground bidirectional
rlabel metal5 s -3283 3773 303275 4083 6 vssd1
port 315 nsew ground bidirectional
rlabel metal5 s -3283 21773 303275 22083 6 vssd1
port 315 nsew ground bidirectional
rlabel metal5 s -3283 39773 303275 40083 6 vssd1
port 315 nsew ground bidirectional
rlabel metal5 s -3283 57773 303275 58083 6 vssd1
port 315 nsew ground bidirectional
rlabel metal5 s -3283 75773 303275 76083 6 vssd1
port 315 nsew ground bidirectional
rlabel metal5 s -3283 93773 303275 94083 6 vssd1
port 315 nsew ground bidirectional
rlabel metal5 s -3283 111773 303275 112083 6 vssd1
port 315 nsew ground bidirectional
rlabel metal5 s -3283 129773 303275 130083 6 vssd1
port 315 nsew ground bidirectional
rlabel metal5 s -3283 147773 303275 148083 6 vssd1
port 315 nsew ground bidirectional
rlabel metal5 s -3283 165773 303275 166083 6 vssd1
port 315 nsew ground bidirectional
rlabel metal5 s -3283 183773 303275 184083 6 vssd1
port 315 nsew ground bidirectional
rlabel metal5 s -3283 201773 303275 202083 6 vssd1
port 315 nsew ground bidirectional
rlabel metal5 s -3283 219773 303275 220083 6 vssd1
port 315 nsew ground bidirectional
rlabel metal5 s -3283 237773 303275 238083 6 vssd1
port 315 nsew ground bidirectional
rlabel metal5 s -3283 255773 303275 256083 6 vssd1
port 315 nsew ground bidirectional
rlabel metal5 s -3283 273773 303275 274083 6 vssd1
port 315 nsew ground bidirectional
rlabel metal5 s -3283 291773 303275 292083 6 vssd1
port 315 nsew ground bidirectional
rlabel metal4 s -2323 -1427 -2013 301307 4 vssd2
port 316 nsew ground bidirectional
rlabel metal5 s -2323 -1427 302315 -1117 8 vssd2
port 316 nsew ground bidirectional
rlabel metal5 s -2323 300997 302315 301307 6 vssd2
port 316 nsew ground bidirectional
rlabel metal4 s 302005 -1427 302315 301307 6 vssd2
port 316 nsew ground bidirectional
rlabel metal4 s 6597 -2387 6907 302267 6 vssd2
port 316 nsew ground bidirectional
rlabel metal4 s 24597 -2387 24907 302267 6 vssd2
port 316 nsew ground bidirectional
rlabel metal4 s 42597 -2387 42907 51721 6 vssd2
port 316 nsew ground bidirectional
rlabel metal4 s 42597 59415 42907 82289 6 vssd2
port 316 nsew ground bidirectional
rlabel metal4 s 42597 94967 42907 302267 6 vssd2
port 316 nsew ground bidirectional
rlabel metal4 s 60597 -2387 60907 302267 6 vssd2
port 316 nsew ground bidirectional
rlabel metal4 s 78597 -2387 78907 302267 6 vssd2
port 316 nsew ground bidirectional
rlabel metal4 s 96597 -2387 96907 302267 6 vssd2
port 316 nsew ground bidirectional
rlabel metal4 s 114597 -2387 114907 302267 6 vssd2
port 316 nsew ground bidirectional
rlabel metal4 s 132597 -2387 132907 302267 6 vssd2
port 316 nsew ground bidirectional
rlabel metal4 s 150597 -2387 150907 302267 6 vssd2
port 316 nsew ground bidirectional
rlabel metal4 s 168597 -2387 168907 302267 6 vssd2
port 316 nsew ground bidirectional
rlabel metal4 s 186597 -2387 186907 302267 6 vssd2
port 316 nsew ground bidirectional
rlabel metal4 s 204597 -2387 204907 302267 6 vssd2
port 316 nsew ground bidirectional
rlabel metal4 s 222597 -2387 222907 302267 6 vssd2
port 316 nsew ground bidirectional
rlabel metal4 s 240597 -2387 240907 302267 6 vssd2
port 316 nsew ground bidirectional
rlabel metal4 s 258597 -2387 258907 302267 6 vssd2
port 316 nsew ground bidirectional
rlabel metal4 s 276597 -2387 276907 302267 6 vssd2
port 316 nsew ground bidirectional
rlabel metal4 s 294597 -2387 294907 302267 6 vssd2
port 316 nsew ground bidirectional
rlabel metal5 s -3283 7493 303275 7803 6 vssd2
port 316 nsew ground bidirectional
rlabel metal5 s -3283 25493 303275 25803 6 vssd2
port 316 nsew ground bidirectional
rlabel metal5 s -3283 43493 303275 43803 6 vssd2
port 316 nsew ground bidirectional
rlabel metal5 s -3283 61493 303275 61803 6 vssd2
port 316 nsew ground bidirectional
rlabel metal5 s -3283 79493 303275 79803 6 vssd2
port 316 nsew ground bidirectional
rlabel metal5 s -3283 97493 303275 97803 6 vssd2
port 316 nsew ground bidirectional
rlabel metal5 s -3283 115493 303275 115803 6 vssd2
port 316 nsew ground bidirectional
rlabel metal5 s -3283 133493 303275 133803 6 vssd2
port 316 nsew ground bidirectional
rlabel metal5 s -3283 151493 303275 151803 6 vssd2
port 316 nsew ground bidirectional
rlabel metal5 s -3283 169493 303275 169803 6 vssd2
port 316 nsew ground bidirectional
rlabel metal5 s -3283 187493 303275 187803 6 vssd2
port 316 nsew ground bidirectional
rlabel metal5 s -3283 205493 303275 205803 6 vssd2
port 316 nsew ground bidirectional
rlabel metal5 s -3283 223493 303275 223803 6 vssd2
port 316 nsew ground bidirectional
rlabel metal5 s -3283 241493 303275 241803 6 vssd2
port 316 nsew ground bidirectional
rlabel metal5 s -3283 259493 303275 259803 6 vssd2
port 316 nsew ground bidirectional
rlabel metal5 s -3283 277493 303275 277803 6 vssd2
port 316 nsew ground bidirectional
rlabel metal5 s -3283 295493 303275 295803 6 vssd2
port 316 nsew ground bidirectional
rlabel metal2 s 11900 -480 12012 240 8 wb_clk_i
port 317 nsew signal input
rlabel metal2 s 12460 -480 12572 240 8 wb_rst_i
port 318 nsew signal input
rlabel metal2 s 13020 -480 13132 240 8 wbs_ack_o
port 319 nsew signal output
rlabel metal2 s 15260 -480 15372 240 8 wbs_adr_i[0]
port 320 nsew signal input
rlabel metal2 s 34300 -480 34412 240 8 wbs_adr_i[10]
port 321 nsew signal input
rlabel metal2 s 35980 -480 36092 240 8 wbs_adr_i[11]
port 322 nsew signal input
rlabel metal2 s 37660 -480 37772 240 8 wbs_adr_i[12]
port 323 nsew signal input
rlabel metal2 s 39340 -480 39452 240 8 wbs_adr_i[13]
port 324 nsew signal input
rlabel metal2 s 41020 -480 41132 240 8 wbs_adr_i[14]
port 325 nsew signal input
rlabel metal2 s 42700 -480 42812 240 8 wbs_adr_i[15]
port 326 nsew signal input
rlabel metal2 s 44380 -480 44492 240 8 wbs_adr_i[16]
port 327 nsew signal input
rlabel metal2 s 46060 -480 46172 240 8 wbs_adr_i[17]
port 328 nsew signal input
rlabel metal2 s 47740 -480 47852 240 8 wbs_adr_i[18]
port 329 nsew signal input
rlabel metal2 s 49420 -480 49532 240 8 wbs_adr_i[19]
port 330 nsew signal input
rlabel metal2 s 17500 -480 17612 240 8 wbs_adr_i[1]
port 331 nsew signal input
rlabel metal2 s 51100 -480 51212 240 8 wbs_adr_i[20]
port 332 nsew signal input
rlabel metal2 s 52780 -480 52892 240 8 wbs_adr_i[21]
port 333 nsew signal input
rlabel metal2 s 54460 -480 54572 240 8 wbs_adr_i[22]
port 334 nsew signal input
rlabel metal2 s 56140 -480 56252 240 8 wbs_adr_i[23]
port 335 nsew signal input
rlabel metal2 s 57820 -480 57932 240 8 wbs_adr_i[24]
port 336 nsew signal input
rlabel metal2 s 59500 -480 59612 240 8 wbs_adr_i[25]
port 337 nsew signal input
rlabel metal2 s 61180 -480 61292 240 8 wbs_adr_i[26]
port 338 nsew signal input
rlabel metal2 s 62860 -480 62972 240 8 wbs_adr_i[27]
port 339 nsew signal input
rlabel metal2 s 64540 -480 64652 240 8 wbs_adr_i[28]
port 340 nsew signal input
rlabel metal2 s 66220 -480 66332 240 8 wbs_adr_i[29]
port 341 nsew signal input
rlabel metal2 s 19740 -480 19852 240 8 wbs_adr_i[2]
port 342 nsew signal input
rlabel metal2 s 67900 -480 68012 240 8 wbs_adr_i[30]
port 343 nsew signal input
rlabel metal2 s 69580 -480 69692 240 8 wbs_adr_i[31]
port 344 nsew signal input
rlabel metal2 s 21980 -480 22092 240 8 wbs_adr_i[3]
port 345 nsew signal input
rlabel metal2 s 24220 -480 24332 240 8 wbs_adr_i[4]
port 346 nsew signal input
rlabel metal2 s 25900 -480 26012 240 8 wbs_adr_i[5]
port 347 nsew signal input
rlabel metal2 s 27580 -480 27692 240 8 wbs_adr_i[6]
port 348 nsew signal input
rlabel metal2 s 29260 -480 29372 240 8 wbs_adr_i[7]
port 349 nsew signal input
rlabel metal2 s 30940 -480 31052 240 8 wbs_adr_i[8]
port 350 nsew signal input
rlabel metal2 s 32620 -480 32732 240 8 wbs_adr_i[9]
port 351 nsew signal input
rlabel metal2 s 13580 -480 13692 240 8 wbs_cyc_i
port 352 nsew signal input
rlabel metal2 s 15820 -480 15932 240 8 wbs_dat_i[0]
port 353 nsew signal input
rlabel metal2 s 34860 -480 34972 240 8 wbs_dat_i[10]
port 354 nsew signal input
rlabel metal2 s 36540 -480 36652 240 8 wbs_dat_i[11]
port 355 nsew signal input
rlabel metal2 s 38220 -480 38332 240 8 wbs_dat_i[12]
port 356 nsew signal input
rlabel metal2 s 39900 -480 40012 240 8 wbs_dat_i[13]
port 357 nsew signal input
rlabel metal2 s 41580 -480 41692 240 8 wbs_dat_i[14]
port 358 nsew signal input
rlabel metal2 s 43260 -480 43372 240 8 wbs_dat_i[15]
port 359 nsew signal input
rlabel metal2 s 44940 -480 45052 240 8 wbs_dat_i[16]
port 360 nsew signal input
rlabel metal2 s 46620 -480 46732 240 8 wbs_dat_i[17]
port 361 nsew signal input
rlabel metal2 s 48300 -480 48412 240 8 wbs_dat_i[18]
port 362 nsew signal input
rlabel metal2 s 49980 -480 50092 240 8 wbs_dat_i[19]
port 363 nsew signal input
rlabel metal2 s 18060 -480 18172 240 8 wbs_dat_i[1]
port 364 nsew signal input
rlabel metal2 s 51660 -480 51772 240 8 wbs_dat_i[20]
port 365 nsew signal input
rlabel metal2 s 53340 -480 53452 240 8 wbs_dat_i[21]
port 366 nsew signal input
rlabel metal2 s 55020 -480 55132 240 8 wbs_dat_i[22]
port 367 nsew signal input
rlabel metal2 s 56700 -480 56812 240 8 wbs_dat_i[23]
port 368 nsew signal input
rlabel metal2 s 58380 -480 58492 240 8 wbs_dat_i[24]
port 369 nsew signal input
rlabel metal2 s 60060 -480 60172 240 8 wbs_dat_i[25]
port 370 nsew signal input
rlabel metal2 s 61740 -480 61852 240 8 wbs_dat_i[26]
port 371 nsew signal input
rlabel metal2 s 63420 -480 63532 240 8 wbs_dat_i[27]
port 372 nsew signal input
rlabel metal2 s 65100 -480 65212 240 8 wbs_dat_i[28]
port 373 nsew signal input
rlabel metal2 s 66780 -480 66892 240 8 wbs_dat_i[29]
port 374 nsew signal input
rlabel metal2 s 20300 -480 20412 240 8 wbs_dat_i[2]
port 375 nsew signal input
rlabel metal2 s 68460 -480 68572 240 8 wbs_dat_i[30]
port 376 nsew signal input
rlabel metal2 s 70140 -480 70252 240 8 wbs_dat_i[31]
port 377 nsew signal input
rlabel metal2 s 22540 -480 22652 240 8 wbs_dat_i[3]
port 378 nsew signal input
rlabel metal2 s 24780 -480 24892 240 8 wbs_dat_i[4]
port 379 nsew signal input
rlabel metal2 s 26460 -480 26572 240 8 wbs_dat_i[5]
port 380 nsew signal input
rlabel metal2 s 28140 -480 28252 240 8 wbs_dat_i[6]
port 381 nsew signal input
rlabel metal2 s 29820 -480 29932 240 8 wbs_dat_i[7]
port 382 nsew signal input
rlabel metal2 s 31500 -480 31612 240 8 wbs_dat_i[8]
port 383 nsew signal input
rlabel metal2 s 33180 -480 33292 240 8 wbs_dat_i[9]
port 384 nsew signal input
rlabel metal2 s 16380 -480 16492 240 8 wbs_dat_o[0]
port 385 nsew signal output
rlabel metal2 s 35420 -480 35532 240 8 wbs_dat_o[10]
port 386 nsew signal output
rlabel metal2 s 37100 -480 37212 240 8 wbs_dat_o[11]
port 387 nsew signal output
rlabel metal2 s 38780 -480 38892 240 8 wbs_dat_o[12]
port 388 nsew signal output
rlabel metal2 s 40460 -480 40572 240 8 wbs_dat_o[13]
port 389 nsew signal output
rlabel metal2 s 42140 -480 42252 240 8 wbs_dat_o[14]
port 390 nsew signal output
rlabel metal2 s 43820 -480 43932 240 8 wbs_dat_o[15]
port 391 nsew signal output
rlabel metal2 s 45500 -480 45612 240 8 wbs_dat_o[16]
port 392 nsew signal output
rlabel metal2 s 47180 -480 47292 240 8 wbs_dat_o[17]
port 393 nsew signal output
rlabel metal2 s 48860 -480 48972 240 8 wbs_dat_o[18]
port 394 nsew signal output
rlabel metal2 s 50540 -480 50652 240 8 wbs_dat_o[19]
port 395 nsew signal output
rlabel metal2 s 18620 -480 18732 240 8 wbs_dat_o[1]
port 396 nsew signal output
rlabel metal2 s 52220 -480 52332 240 8 wbs_dat_o[20]
port 397 nsew signal output
rlabel metal2 s 53900 -480 54012 240 8 wbs_dat_o[21]
port 398 nsew signal output
rlabel metal2 s 55580 -480 55692 240 8 wbs_dat_o[22]
port 399 nsew signal output
rlabel metal2 s 57260 -480 57372 240 8 wbs_dat_o[23]
port 400 nsew signal output
rlabel metal2 s 58940 -480 59052 240 8 wbs_dat_o[24]
port 401 nsew signal output
rlabel metal2 s 60620 -480 60732 240 8 wbs_dat_o[25]
port 402 nsew signal output
rlabel metal2 s 62300 -480 62412 240 8 wbs_dat_o[26]
port 403 nsew signal output
rlabel metal2 s 63980 -480 64092 240 8 wbs_dat_o[27]
port 404 nsew signal output
rlabel metal2 s 65660 -480 65772 240 8 wbs_dat_o[28]
port 405 nsew signal output
rlabel metal2 s 67340 -480 67452 240 8 wbs_dat_o[29]
port 406 nsew signal output
rlabel metal2 s 20860 -480 20972 240 8 wbs_dat_o[2]
port 407 nsew signal output
rlabel metal2 s 69020 -480 69132 240 8 wbs_dat_o[30]
port 408 nsew signal output
rlabel metal2 s 70700 -480 70812 240 8 wbs_dat_o[31]
port 409 nsew signal output
rlabel metal2 s 23100 -480 23212 240 8 wbs_dat_o[3]
port 410 nsew signal output
rlabel metal2 s 25340 -480 25452 240 8 wbs_dat_o[4]
port 411 nsew signal output
rlabel metal2 s 27020 -480 27132 240 8 wbs_dat_o[5]
port 412 nsew signal output
rlabel metal2 s 28700 -480 28812 240 8 wbs_dat_o[6]
port 413 nsew signal output
rlabel metal2 s 30380 -480 30492 240 8 wbs_dat_o[7]
port 414 nsew signal output
rlabel metal2 s 32060 -480 32172 240 8 wbs_dat_o[8]
port 415 nsew signal output
rlabel metal2 s 33740 -480 33852 240 8 wbs_dat_o[9]
port 416 nsew signal output
rlabel metal2 s 16940 -480 17052 240 8 wbs_sel_i[0]
port 417 nsew signal input
rlabel metal2 s 19180 -480 19292 240 8 wbs_sel_i[1]
port 418 nsew signal input
rlabel metal2 s 21420 -480 21532 240 8 wbs_sel_i[2]
port 419 nsew signal input
rlabel metal2 s 23660 -480 23772 240 8 wbs_sel_i[3]
port 420 nsew signal input
rlabel metal2 s 14140 -480 14252 240 8 wbs_stb_i
port 421 nsew signal input
rlabel metal2 s 14700 -480 14812 240 8 wbs_we_i
port 422 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 300000 300000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 6858984
string GDS_FILE /home/maltik/uP16_gfmpw/openlane/user_project_wrapper/runs/22_12_05_08_36/results/signoff/user_project_wrapper.magic.gds
string GDS_START 4105142
<< end >>

